module sinusoid_ROM (
  input               clk,
  input      [11:0] raddr,
  output     [23:0]  dout
  );
 
 //ROM memory storing 4096 samples addressable
 //on 12 bit address (raddr)
reg signed [23:0] sine_sample;

always @(posedge clk)
begin
case(raddr)
 0: sine_sample <= 0;
 1: sine_sample <= 1609;
 2: sine_sample <= 3217;
 3: sine_sample <= 4826;
 4: sine_sample <= 6434;
 5: sine_sample <= 8043;
 6: sine_sample <= 9651;
 7: sine_sample <= 11259;
 8: sine_sample <= 12868;
 9: sine_sample <= 14476;
 10: sine_sample <= 16084;
 11: sine_sample <= 17693;
 12: sine_sample <= 19301;
 13: sine_sample <= 20909;
 14: sine_sample <= 22517;
 15: sine_sample <= 24125;
 16: sine_sample <= 25733;
 17: sine_sample <= 27341;
 18: sine_sample <= 28949;
 19: sine_sample <= 30557;
 20: sine_sample <= 32165;
 21: sine_sample <= 33773;
 22: sine_sample <= 35380;
 23: sine_sample <= 36988;
 24: sine_sample <= 38595;
 25: sine_sample <= 40203;
 26: sine_sample <= 41810;
 27: sine_sample <= 43417;
 28: sine_sample <= 45024;
 29: sine_sample <= 46631;
 30: sine_sample <= 48238;
 31: sine_sample <= 49845;
 32: sine_sample <= 51451;
 33: sine_sample <= 53058;
 34: sine_sample <= 54664;
 35: sine_sample <= 56270;
 36: sine_sample <= 57877;
 37: sine_sample <= 59483;
 38: sine_sample <= 61088;
 39: sine_sample <= 62694;
 40: sine_sample <= 64300;
 41: sine_sample <= 65905;
 42: sine_sample <= 67510;
 43: sine_sample <= 69115;
 44: sine_sample <= 70720;
 45: sine_sample <= 72325;
 46: sine_sample <= 73930;
 47: sine_sample <= 75534;
 48: sine_sample <= 77138;
 49: sine_sample <= 78742;
 50: sine_sample <= 80346;
 51: sine_sample <= 81950;
 52: sine_sample <= 83553;
 53: sine_sample <= 85156;
 54: sine_sample <= 86760;
 55: sine_sample <= 88362;
 56: sine_sample <= 89965;
 57: sine_sample <= 91568;
 58: sine_sample <= 93170;
 59: sine_sample <= 94772;
 60: sine_sample <= 96374;
 61: sine_sample <= 97975;
 62: sine_sample <= 99577;
 63: sine_sample <= 101178;
 64: sine_sample <= 102779;
 65: sine_sample <= 104379;
 66: sine_sample <= 105980;
 67: sine_sample <= 107580;
 68: sine_sample <= 109180;
 69: sine_sample <= 110779;
 70: sine_sample <= 112379;
 71: sine_sample <= 113978;
 72: sine_sample <= 115576;
 73: sine_sample <= 117175;
 74: sine_sample <= 118773;
 75: sine_sample <= 120371;
 76: sine_sample <= 121969;
 77: sine_sample <= 123566;
 78: sine_sample <= 125164;
 79: sine_sample <= 126760;
 80: sine_sample <= 128357;
 81: sine_sample <= 129953;
 82: sine_sample <= 131549;
 83: sine_sample <= 133145;
 84: sine_sample <= 134740;
 85: sine_sample <= 136335;
 86: sine_sample <= 137930;
 87: sine_sample <= 139524;
 88: sine_sample <= 141118;
 89: sine_sample <= 142712;
 90: sine_sample <= 144305;
 91: sine_sample <= 145898;
 92: sine_sample <= 147491;
 93: sine_sample <= 149083;
 94: sine_sample <= 150675;
 95: sine_sample <= 152267;
 96: sine_sample <= 153858;
 97: sine_sample <= 155449;
 98: sine_sample <= 157040;
 99: sine_sample <= 158630;
 100: sine_sample <= 160220;
 101: sine_sample <= 161809;
 102: sine_sample <= 163398;
 103: sine_sample <= 164987;
 104: sine_sample <= 166575;
 105: sine_sample <= 168163;
 106: sine_sample <= 169750;
 107: sine_sample <= 171337;
 108: sine_sample <= 172924;
 109: sine_sample <= 174510;
 110: sine_sample <= 176096;
 111: sine_sample <= 177682;
 112: sine_sample <= 179267;
 113: sine_sample <= 180851;
 114: sine_sample <= 182435;
 115: sine_sample <= 184019;
 116: sine_sample <= 185603;
 117: sine_sample <= 187185;
 118: sine_sample <= 188768;
 119: sine_sample <= 190350;
 120: sine_sample <= 191931;
 121: sine_sample <= 193512;
 122: sine_sample <= 195093;
 123: sine_sample <= 196673;
 124: sine_sample <= 198253;
 125: sine_sample <= 199832;
 126: sine_sample <= 201411;
 127: sine_sample <= 202989;
 128: sine_sample <= 204567;
 129: sine_sample <= 206145;
 130: sine_sample <= 207721;
 131: sine_sample <= 209298;
 132: sine_sample <= 210874;
 133: sine_sample <= 212449;
 134: sine_sample <= 214024;
 135: sine_sample <= 215598;
 136: sine_sample <= 217172;
 137: sine_sample <= 218746;
 138: sine_sample <= 220318;
 139: sine_sample <= 221891;
 140: sine_sample <= 223462;
 141: sine_sample <= 225034;
 142: sine_sample <= 226605;
 143: sine_sample <= 228175;
 144: sine_sample <= 229744;
 145: sine_sample <= 231314;
 146: sine_sample <= 232882;
 147: sine_sample <= 234450;
 148: sine_sample <= 236018;
 149: sine_sample <= 237585;
 150: sine_sample <= 239151;
 151: sine_sample <= 240717;
 152: sine_sample <= 242282;
 153: sine_sample <= 243847;
 154: sine_sample <= 245411;
 155: sine_sample <= 246974;
 156: sine_sample <= 248537;
 157: sine_sample <= 250100;
 158: sine_sample <= 251662;
 159: sine_sample <= 253223;
 160: sine_sample <= 254783;
 161: sine_sample <= 256343;
 162: sine_sample <= 257903;
 163: sine_sample <= 259461;
 164: sine_sample <= 261020;
 165: sine_sample <= 262577;
 166: sine_sample <= 264134;
 167: sine_sample <= 265690;
 168: sine_sample <= 267246;
 169: sine_sample <= 268801;
 170: sine_sample <= 270356;
 171: sine_sample <= 271909;
 172: sine_sample <= 273463;
 173: sine_sample <= 275015;
 174: sine_sample <= 276567;
 175: sine_sample <= 278118;
 176: sine_sample <= 279669;
 177: sine_sample <= 281219;
 178: sine_sample <= 282768;
 179: sine_sample <= 284316;
 180: sine_sample <= 285864;
 181: sine_sample <= 287412;
 182: sine_sample <= 288958;
 183: sine_sample <= 290504;
 184: sine_sample <= 292049;
 185: sine_sample <= 293594;
 186: sine_sample <= 295138;
 187: sine_sample <= 296681;
 188: sine_sample <= 298223;
 189: sine_sample <= 299765;
 190: sine_sample <= 301306;
 191: sine_sample <= 302846;
 192: sine_sample <= 304386;
 193: sine_sample <= 305925;
 194: sine_sample <= 307463;
 195: sine_sample <= 309000;
 196: sine_sample <= 310537;
 197: sine_sample <= 312073;
 198: sine_sample <= 313608;
 199: sine_sample <= 315143;
 200: sine_sample <= 316676;
 201: sine_sample <= 318209;
 202: sine_sample <= 319742;
 203: sine_sample <= 321273;
 204: sine_sample <= 322804;
 205: sine_sample <= 324334;
 206: sine_sample <= 325863;
 207: sine_sample <= 327392;
 208: sine_sample <= 328919;
 209: sine_sample <= 330446;
 210: sine_sample <= 331972;
 211: sine_sample <= 333498;
 212: sine_sample <= 335022;
 213: sine_sample <= 336546;
 214: sine_sample <= 338069;
 215: sine_sample <= 339591;
 216: sine_sample <= 341113;
 217: sine_sample <= 342633;
 218: sine_sample <= 344153;
 219: sine_sample <= 345672;
 220: sine_sample <= 347190;
 221: sine_sample <= 348708;
 222: sine_sample <= 350224;
 223: sine_sample <= 351740;
 224: sine_sample <= 353255;
 225: sine_sample <= 354769;
 226: sine_sample <= 356282;
 227: sine_sample <= 357794;
 228: sine_sample <= 359306;
 229: sine_sample <= 360817;
 230: sine_sample <= 362326;
 231: sine_sample <= 363835;
 232: sine_sample <= 365344;
 233: sine_sample <= 366851;
 234: sine_sample <= 368357;
 235: sine_sample <= 369863;
 236: sine_sample <= 371367;
 237: sine_sample <= 372871;
 238: sine_sample <= 374374;
 239: sine_sample <= 375876;
 240: sine_sample <= 377377;
 241: sine_sample <= 378878;
 242: sine_sample <= 380377;
 243: sine_sample <= 381876;
 244: sine_sample <= 383373;
 245: sine_sample <= 384870;
 246: sine_sample <= 386366;
 247: sine_sample <= 387860;
 248: sine_sample <= 389354;
 249: sine_sample <= 390847;
 250: sine_sample <= 392340;
 251: sine_sample <= 393831;
 252: sine_sample <= 395321;
 253: sine_sample <= 396810;
 254: sine_sample <= 398299;
 255: sine_sample <= 399786;
 256: sine_sample <= 401273;
 257: sine_sample <= 402758;
 258: sine_sample <= 404243;
 259: sine_sample <= 405727;
 260: sine_sample <= 407209;
 261: sine_sample <= 408691;
 262: sine_sample <= 410172;
 263: sine_sample <= 411652;
 264: sine_sample <= 413131;
 265: sine_sample <= 414609;
 266: sine_sample <= 416086;
 267: sine_sample <= 417562;
 268: sine_sample <= 419036;
 269: sine_sample <= 420510;
 270: sine_sample <= 421983;
 271: sine_sample <= 423455;
 272: sine_sample <= 424926;
 273: sine_sample <= 426396;
 274: sine_sample <= 427865;
 275: sine_sample <= 429333;
 276: sine_sample <= 430800;
 277: sine_sample <= 432266;
 278: sine_sample <= 433731;
 279: sine_sample <= 435195;
 280: sine_sample <= 436658;
 281: sine_sample <= 438120;
 282: sine_sample <= 439581;
 283: sine_sample <= 441041;
 284: sine_sample <= 442499;
 285: sine_sample <= 443957;
 286: sine_sample <= 445414;
 287: sine_sample <= 446870;
 288: sine_sample <= 448324;
 289: sine_sample <= 449778;
 290: sine_sample <= 451230;
 291: sine_sample <= 452682;
 292: sine_sample <= 454132;
 293: sine_sample <= 455581;
 294: sine_sample <= 457029;
 295: sine_sample <= 458477;
 296: sine_sample <= 459923;
 297: sine_sample <= 461368;
 298: sine_sample <= 462811;
 299: sine_sample <= 464254;
 300: sine_sample <= 465696;
 301: sine_sample <= 467137;
 302: sine_sample <= 468576;
 303: sine_sample <= 470014;
 304: sine_sample <= 471452;
 305: sine_sample <= 472888;
 306: sine_sample <= 474323;
 307: sine_sample <= 475757;
 308: sine_sample <= 477190;
 309: sine_sample <= 478622;
 310: sine_sample <= 480052;
 311: sine_sample <= 481482;
 312: sine_sample <= 482910;
 313: sine_sample <= 484337;
 314: sine_sample <= 485763;
 315: sine_sample <= 487188;
 316: sine_sample <= 488612;
 317: sine_sample <= 490035;
 318: sine_sample <= 491456;
 319: sine_sample <= 492876;
 320: sine_sample <= 494295;
 321: sine_sample <= 495713;
 322: sine_sample <= 497130;
 323: sine_sample <= 498546;
 324: sine_sample <= 499960;
 325: sine_sample <= 501374;
 326: sine_sample <= 502786;
 327: sine_sample <= 504197;
 328: sine_sample <= 505606;
 329: sine_sample <= 507015;
 330: sine_sample <= 508422;
 331: sine_sample <= 509829;
 332: sine_sample <= 511234;
 333: sine_sample <= 512637;
 334: sine_sample <= 514040;
 335: sine_sample <= 515441;
 336: sine_sample <= 516841;
 337: sine_sample <= 518240;
 338: sine_sample <= 519638;
 339: sine_sample <= 521034;
 340: sine_sample <= 522430;
 341: sine_sample <= 523824;
 342: sine_sample <= 525217;
 343: sine_sample <= 526608;
 344: sine_sample <= 527998;
 345: sine_sample <= 529387;
 346: sine_sample <= 530775;
 347: sine_sample <= 532162;
 348: sine_sample <= 533547;
 349: sine_sample <= 534931;
 350: sine_sample <= 536314;
 351: sine_sample <= 537696;
 352: sine_sample <= 539076;
 353: sine_sample <= 540455;
 354: sine_sample <= 541833;
 355: sine_sample <= 543209;
 356: sine_sample <= 544584;
 357: sine_sample <= 545958;
 358: sine_sample <= 547331;
 359: sine_sample <= 548702;
 360: sine_sample <= 550072;
 361: sine_sample <= 551441;
 362: sine_sample <= 552808;
 363: sine_sample <= 554175;
 364: sine_sample <= 555539;
 365: sine_sample <= 556903;
 366: sine_sample <= 558265;
 367: sine_sample <= 559626;
 368: sine_sample <= 560986;
 369: sine_sample <= 562344;
 370: sine_sample <= 563701;
 371: sine_sample <= 565057;
 372: sine_sample <= 566411;
 373: sine_sample <= 567764;
 374: sine_sample <= 569116;
 375: sine_sample <= 570466;
 376: sine_sample <= 571815;
 377: sine_sample <= 573162;
 378: sine_sample <= 574509;
 379: sine_sample <= 575854;
 380: sine_sample <= 577197;
 381: sine_sample <= 578539;
 382: sine_sample <= 579880;
 383: sine_sample <= 581220;
 384: sine_sample <= 582558;
 385: sine_sample <= 583894;
 386: sine_sample <= 585230;
 387: sine_sample <= 586564;
 388: sine_sample <= 587896;
 389: sine_sample <= 589228;
 390: sine_sample <= 590557;
 391: sine_sample <= 591886;
 392: sine_sample <= 593213;
 393: sine_sample <= 594539;
 394: sine_sample <= 595863;
 395: sine_sample <= 597186;
 396: sine_sample <= 598507;
 397: sine_sample <= 599827;
 398: sine_sample <= 601146;
 399: sine_sample <= 602463;
 400: sine_sample <= 603779;
 401: sine_sample <= 605093;
 402: sine_sample <= 606406;
 403: sine_sample <= 607718;
 404: sine_sample <= 609028;
 405: sine_sample <= 610336;
 406: sine_sample <= 611644;
 407: sine_sample <= 612949;
 408: sine_sample <= 614254;
 409: sine_sample <= 615557;
 410: sine_sample <= 616858;
 411: sine_sample <= 618158;
 412: sine_sample <= 619457;
 413: sine_sample <= 620754;
 414: sine_sample <= 622049;
 415: sine_sample <= 623343;
 416: sine_sample <= 624636;
 417: sine_sample <= 625927;
 418: sine_sample <= 627217;
 419: sine_sample <= 628505;
 420: sine_sample <= 629792;
 421: sine_sample <= 631077;
 422: sine_sample <= 632361;
 423: sine_sample <= 633644;
 424: sine_sample <= 634924;
 425: sine_sample <= 636204;
 426: sine_sample <= 637482;
 427: sine_sample <= 638758;
 428: sine_sample <= 640033;
 429: sine_sample <= 641306;
 430: sine_sample <= 642578;
 431: sine_sample <= 643848;
 432: sine_sample <= 645117;
 433: sine_sample <= 646384;
 434: sine_sample <= 647650;
 435: sine_sample <= 648915;
 436: sine_sample <= 650177;
 437: sine_sample <= 651438;
 438: sine_sample <= 652698;
 439: sine_sample <= 653956;
 440: sine_sample <= 655213;
 441: sine_sample <= 656468;
 442: sine_sample <= 657721;
 443: sine_sample <= 658973;
 444: sine_sample <= 660224;
 445: sine_sample <= 661473;
 446: sine_sample <= 662720;
 447: sine_sample <= 663966;
 448: sine_sample <= 665210;
 449: sine_sample <= 666452;
 450: sine_sample <= 667693;
 451: sine_sample <= 668933;
 452: sine_sample <= 670171;
 453: sine_sample <= 671407;
 454: sine_sample <= 672642;
 455: sine_sample <= 673875;
 456: sine_sample <= 675106;
 457: sine_sample <= 676336;
 458: sine_sample <= 677565;
 459: sine_sample <= 678792;
 460: sine_sample <= 680017;
 461: sine_sample <= 681240;
 462: sine_sample <= 682462;
 463: sine_sample <= 683683;
 464: sine_sample <= 684901;
 465: sine_sample <= 686119;
 466: sine_sample <= 687334;
 467: sine_sample <= 688548;
 468: sine_sample <= 689760;
 469: sine_sample <= 690971;
 470: sine_sample <= 692180;
 471: sine_sample <= 693388;
 472: sine_sample <= 694593;
 473: sine_sample <= 695798;
 474: sine_sample <= 697000;
 475: sine_sample <= 698201;
 476: sine_sample <= 699400;
 477: sine_sample <= 700598;
 478: sine_sample <= 701794;
 479: sine_sample <= 702988;
 480: sine_sample <= 704181;
 481: sine_sample <= 705372;
 482: sine_sample <= 706561;
 483: sine_sample <= 707749;
 484: sine_sample <= 708935;
 485: sine_sample <= 710119;
 486: sine_sample <= 711302;
 487: sine_sample <= 712483;
 488: sine_sample <= 713662;
 489: sine_sample <= 714840;
 490: sine_sample <= 716016;
 491: sine_sample <= 717190;
 492: sine_sample <= 718362;
 493: sine_sample <= 719533;
 494: sine_sample <= 720702;
 495: sine_sample <= 721870;
 496: sine_sample <= 723036;
 497: sine_sample <= 724200;
 498: sine_sample <= 725362;
 499: sine_sample <= 726523;
 500: sine_sample <= 727682;
 501: sine_sample <= 728839;
 502: sine_sample <= 729995;
 503: sine_sample <= 731149;
 504: sine_sample <= 732301;
 505: sine_sample <= 733451;
 506: sine_sample <= 734600;
 507: sine_sample <= 735747;
 508: sine_sample <= 736892;
 509: sine_sample <= 738035;
 510: sine_sample <= 739177;
 511: sine_sample <= 740317;
 512: sine_sample <= 741455;
 513: sine_sample <= 742592;
 514: sine_sample <= 743727;
 515: sine_sample <= 744860;
 516: sine_sample <= 745991;
 517: sine_sample <= 747120;
 518: sine_sample <= 748248;
 519: sine_sample <= 749374;
 520: sine_sample <= 750498;
 521: sine_sample <= 751621;
 522: sine_sample <= 752741;
 523: sine_sample <= 753860;
 524: sine_sample <= 754977;
 525: sine_sample <= 756093;
 526: sine_sample <= 757206;
 527: sine_sample <= 758318;
 528: sine_sample <= 759428;
 529: sine_sample <= 760536;
 530: sine_sample <= 761643;
 531: sine_sample <= 762748;
 532: sine_sample <= 763850;
 533: sine_sample <= 764951;
 534: sine_sample <= 766051;
 535: sine_sample <= 767148;
 536: sine_sample <= 768244;
 537: sine_sample <= 769338;
 538: sine_sample <= 770430;
 539: sine_sample <= 771520;
 540: sine_sample <= 772608;
 541: sine_sample <= 773695;
 542: sine_sample <= 774780;
 543: sine_sample <= 775863;
 544: sine_sample <= 776944;
 545: sine_sample <= 778023;
 546: sine_sample <= 779100;
 547: sine_sample <= 780176;
 548: sine_sample <= 781250;
 549: sine_sample <= 782322;
 550: sine_sample <= 783392;
 551: sine_sample <= 784460;
 552: sine_sample <= 785527;
 553: sine_sample <= 786591;
 554: sine_sample <= 787654;
 555: sine_sample <= 788715;
 556: sine_sample <= 789774;
 557: sine_sample <= 790831;
 558: sine_sample <= 791886;
 559: sine_sample <= 792940;
 560: sine_sample <= 793991;
 561: sine_sample <= 795041;
 562: sine_sample <= 796089;
 563: sine_sample <= 797135;
 564: sine_sample <= 798179;
 565: sine_sample <= 799221;
 566: sine_sample <= 800261;
 567: sine_sample <= 801300;
 568: sine_sample <= 802336;
 569: sine_sample <= 803371;
 570: sine_sample <= 804404;
 571: sine_sample <= 805434;
 572: sine_sample <= 806463;
 573: sine_sample <= 807491;
 574: sine_sample <= 808516;
 575: sine_sample <= 809539;
 576: sine_sample <= 810560;
 577: sine_sample <= 811580;
 578: sine_sample <= 812597;
 579: sine_sample <= 813613;
 580: sine_sample <= 814627;
 581: sine_sample <= 815639;
 582: sine_sample <= 816648;
 583: sine_sample <= 817656;
 584: sine_sample <= 818662;
 585: sine_sample <= 819667;
 586: sine_sample <= 820669;
 587: sine_sample <= 821669;
 588: sine_sample <= 822667;
 589: sine_sample <= 823664;
 590: sine_sample <= 824658;
 591: sine_sample <= 825651;
 592: sine_sample <= 826641;
 593: sine_sample <= 827630;
 594: sine_sample <= 828617;
 595: sine_sample <= 829601;
 596: sine_sample <= 830584;
 597: sine_sample <= 831565;
 598: sine_sample <= 832544;
 599: sine_sample <= 833521;
 600: sine_sample <= 834496;
 601: sine_sample <= 835469;
 602: sine_sample <= 836440;
 603: sine_sample <= 837409;
 604: sine_sample <= 838376;
 605: sine_sample <= 839341;
 606: sine_sample <= 840304;
 607: sine_sample <= 841265;
 608: sine_sample <= 842224;
 609: sine_sample <= 843181;
 610: sine_sample <= 844137;
 611: sine_sample <= 845090;
 612: sine_sample <= 846041;
 613: sine_sample <= 846990;
 614: sine_sample <= 847938;
 615: sine_sample <= 848883;
 616: sine_sample <= 849826;
 617: sine_sample <= 850767;
 618: sine_sample <= 851707;
 619: sine_sample <= 852644;
 620: sine_sample <= 853579;
 621: sine_sample <= 854512;
 622: sine_sample <= 855444;
 623: sine_sample <= 856373;
 624: sine_sample <= 857300;
 625: sine_sample <= 858225;
 626: sine_sample <= 859148;
 627: sine_sample <= 860069;
 628: sine_sample <= 860989;
 629: sine_sample <= 861906;
 630: sine_sample <= 862821;
 631: sine_sample <= 863734;
 632: sine_sample <= 864645;
 633: sine_sample <= 865554;
 634: sine_sample <= 866461;
 635: sine_sample <= 867365;
 636: sine_sample <= 868268;
 637: sine_sample <= 869169;
 638: sine_sample <= 870068;
 639: sine_sample <= 870965;
 640: sine_sample <= 871859;
 641: sine_sample <= 872752;
 642: sine_sample <= 873642;
 643: sine_sample <= 874531;
 644: sine_sample <= 875417;
 645: sine_sample <= 876302;
 646: sine_sample <= 877184;
 647: sine_sample <= 878064;
 648: sine_sample <= 878942;
 649: sine_sample <= 879819;
 650: sine_sample <= 880693;
 651: sine_sample <= 881565;
 652: sine_sample <= 882434;
 653: sine_sample <= 883302;
 654: sine_sample <= 884168;
 655: sine_sample <= 885032;
 656: sine_sample <= 885893;
 657: sine_sample <= 886753;
 658: sine_sample <= 887610;
 659: sine_sample <= 888466;
 660: sine_sample <= 889319;
 661: sine_sample <= 890170;
 662: sine_sample <= 891019;
 663: sine_sample <= 891866;
 664: sine_sample <= 892711;
 665: sine_sample <= 893553;
 666: sine_sample <= 894394;
 667: sine_sample <= 895233;
 668: sine_sample <= 896069;
 669: sine_sample <= 896903;
 670: sine_sample <= 897736;
 671: sine_sample <= 898566;
 672: sine_sample <= 899394;
 673: sine_sample <= 900220;
 674: sine_sample <= 901043;
 675: sine_sample <= 901865;
 676: sine_sample <= 902685;
 677: sine_sample <= 903502;
 678: sine_sample <= 904317;
 679: sine_sample <= 905130;
 680: sine_sample <= 905941;
 681: sine_sample <= 906750;
 682: sine_sample <= 907557;
 683: sine_sample <= 908362;
 684: sine_sample <= 909164;
 685: sine_sample <= 909964;
 686: sine_sample <= 910763;
 687: sine_sample <= 911559;
 688: sine_sample <= 912352;
 689: sine_sample <= 913144;
 690: sine_sample <= 913934;
 691: sine_sample <= 914721;
 692: sine_sample <= 915507;
 693: sine_sample <= 916290;
 694: sine_sample <= 917071;
 695: sine_sample <= 917850;
 696: sine_sample <= 918626;
 697: sine_sample <= 919401;
 698: sine_sample <= 920173;
 699: sine_sample <= 920943;
 700: sine_sample <= 921711;
 701: sine_sample <= 922477;
 702: sine_sample <= 923241;
 703: sine_sample <= 924002;
 704: sine_sample <= 924762;
 705: sine_sample <= 925519;
 706: sine_sample <= 926274;
 707: sine_sample <= 927027;
 708: sine_sample <= 927777;
 709: sine_sample <= 928526;
 710: sine_sample <= 929272;
 711: sine_sample <= 930016;
 712: sine_sample <= 930758;
 713: sine_sample <= 931497;
 714: sine_sample <= 932235;
 715: sine_sample <= 932970;
 716: sine_sample <= 933703;
 717: sine_sample <= 934434;
 718: sine_sample <= 935163;
 719: sine_sample <= 935889;
 720: sine_sample <= 936614;
 721: sine_sample <= 937336;
 722: sine_sample <= 938056;
 723: sine_sample <= 938773;
 724: sine_sample <= 939489;
 725: sine_sample <= 940202;
 726: sine_sample <= 940913;
 727: sine_sample <= 941622;
 728: sine_sample <= 942329;
 729: sine_sample <= 943033;
 730: sine_sample <= 943735;
 731: sine_sample <= 944435;
 732: sine_sample <= 945133;
 733: sine_sample <= 945828;
 734: sine_sample <= 946522;
 735: sine_sample <= 947213;
 736: sine_sample <= 947902;
 737: sine_sample <= 948588;
 738: sine_sample <= 949273;
 739: sine_sample <= 949955;
 740: sine_sample <= 950635;
 741: sine_sample <= 951312;
 742: sine_sample <= 951988;
 743: sine_sample <= 952661;
 744: sine_sample <= 953332;
 745: sine_sample <= 954001;
 746: sine_sample <= 954667;
 747: sine_sample <= 955331;
 748: sine_sample <= 955993;
 749: sine_sample <= 956653;
 750: sine_sample <= 957310;
 751: sine_sample <= 957966;
 752: sine_sample <= 958619;
 753: sine_sample <= 959269;
 754: sine_sample <= 959918;
 755: sine_sample <= 960564;
 756: sine_sample <= 961208;
 757: sine_sample <= 961849;
 758: sine_sample <= 962489;
 759: sine_sample <= 963126;
 760: sine_sample <= 963761;
 761: sine_sample <= 964393;
 762: sine_sample <= 965024;
 763: sine_sample <= 965652;
 764: sine_sample <= 966278;
 765: sine_sample <= 966901;
 766: sine_sample <= 967522;
 767: sine_sample <= 968141;
 768: sine_sample <= 968758;
 769: sine_sample <= 969372;
 770: sine_sample <= 969985;
 771: sine_sample <= 970594;
 772: sine_sample <= 971202;
 773: sine_sample <= 971807;
 774: sine_sample <= 972410;
 775: sine_sample <= 973011;
 776: sine_sample <= 973609;
 777: sine_sample <= 974205;
 778: sine_sample <= 974799;
 779: sine_sample <= 975391;
 780: sine_sample <= 975980;
 781: sine_sample <= 976567;
 782: sine_sample <= 977152;
 783: sine_sample <= 977734;
 784: sine_sample <= 978314;
 785: sine_sample <= 978892;
 786: sine_sample <= 979467;
 787: sine_sample <= 980040;
 788: sine_sample <= 980611;
 789: sine_sample <= 981180;
 790: sine_sample <= 981746;
 791: sine_sample <= 982310;
 792: sine_sample <= 982871;
 793: sine_sample <= 983431;
 794: sine_sample <= 983988;
 795: sine_sample <= 984542;
 796: sine_sample <= 985095;
 797: sine_sample <= 985645;
 798: sine_sample <= 986192;
 799: sine_sample <= 986738;
 800: sine_sample <= 987281;
 801: sine_sample <= 987821;
 802: sine_sample <= 988360;
 803: sine_sample <= 988896;
 804: sine_sample <= 989430;
 805: sine_sample <= 989961;
 806: sine_sample <= 990490;
 807: sine_sample <= 991017;
 808: sine_sample <= 991541;
 809: sine_sample <= 992063;
 810: sine_sample <= 992583;
 811: sine_sample <= 993101;
 812: sine_sample <= 993616;
 813: sine_sample <= 994128;
 814: sine_sample <= 994639;
 815: sine_sample <= 995147;
 816: sine_sample <= 995653;
 817: sine_sample <= 996156;
 818: sine_sample <= 996657;
 819: sine_sample <= 997156;
 820: sine_sample <= 997652;
 821: sine_sample <= 998146;
 822: sine_sample <= 998638;
 823: sine_sample <= 999127;
 824: sine_sample <= 999614;
 825: sine_sample <= 1000099;
 826: sine_sample <= 1000581;
 827: sine_sample <= 1001061;
 828: sine_sample <= 1001538;
 829: sine_sample <= 1002013;
 830: sine_sample <= 1002486;
 831: sine_sample <= 1002957;
 832: sine_sample <= 1003425;
 833: sine_sample <= 1003891;
 834: sine_sample <= 1004354;
 835: sine_sample <= 1004815;
 836: sine_sample <= 1005274;
 837: sine_sample <= 1005730;
 838: sine_sample <= 1006184;
 839: sine_sample <= 1006635;
 840: sine_sample <= 1007085;
 841: sine_sample <= 1007531;
 842: sine_sample <= 1007976;
 843: sine_sample <= 1008418;
 844: sine_sample <= 1008858;
 845: sine_sample <= 1009295;
 846: sine_sample <= 1009730;
 847: sine_sample <= 1010162;
 848: sine_sample <= 1010593;
 849: sine_sample <= 1011020;
 850: sine_sample <= 1011446;
 851: sine_sample <= 1011869;
 852: sine_sample <= 1012290;
 853: sine_sample <= 1012708;
 854: sine_sample <= 1013124;
 855: sine_sample <= 1013537;
 856: sine_sample <= 1013948;
 857: sine_sample <= 1014357;
 858: sine_sample <= 1014764;
 859: sine_sample <= 1015168;
 860: sine_sample <= 1015569;
 861: sine_sample <= 1015968;
 862: sine_sample <= 1016365;
 863: sine_sample <= 1016760;
 864: sine_sample <= 1017152;
 865: sine_sample <= 1017541;
 866: sine_sample <= 1017928;
 867: sine_sample <= 1018313;
 868: sine_sample <= 1018696;
 869: sine_sample <= 1019076;
 870: sine_sample <= 1019453;
 871: sine_sample <= 1019829;
 872: sine_sample <= 1020202;
 873: sine_sample <= 1020572;
 874: sine_sample <= 1020940;
 875: sine_sample <= 1021306;
 876: sine_sample <= 1021669;
 877: sine_sample <= 1022030;
 878: sine_sample <= 1022388;
 879: sine_sample <= 1022744;
 880: sine_sample <= 1023098;
 881: sine_sample <= 1023449;
 882: sine_sample <= 1023798;
 883: sine_sample <= 1024144;
 884: sine_sample <= 1024488;
 885: sine_sample <= 1024830;
 886: sine_sample <= 1025169;
 887: sine_sample <= 1025506;
 888: sine_sample <= 1025840;
 889: sine_sample <= 1026172;
 890: sine_sample <= 1026502;
 891: sine_sample <= 1026829;
 892: sine_sample <= 1027153;
 893: sine_sample <= 1027476;
 894: sine_sample <= 1027796;
 895: sine_sample <= 1028113;
 896: sine_sample <= 1028428;
 897: sine_sample <= 1028741;
 898: sine_sample <= 1029051;
 899: sine_sample <= 1029359;
 900: sine_sample <= 1029664;
 901: sine_sample <= 1029967;
 902: sine_sample <= 1030267;
 903: sine_sample <= 1030565;
 904: sine_sample <= 1030861;
 905: sine_sample <= 1031154;
 906: sine_sample <= 1031445;
 907: sine_sample <= 1031733;
 908: sine_sample <= 1032019;
 909: sine_sample <= 1032303;
 910: sine_sample <= 1032584;
 911: sine_sample <= 1032862;
 912: sine_sample <= 1033139;
 913: sine_sample <= 1033412;
 914: sine_sample <= 1033684;
 915: sine_sample <= 1033953;
 916: sine_sample <= 1034219;
 917: sine_sample <= 1034483;
 918: sine_sample <= 1034745;
 919: sine_sample <= 1035004;
 920: sine_sample <= 1035261;
 921: sine_sample <= 1035515;
 922: sine_sample <= 1035767;
 923: sine_sample <= 1036016;
 924: sine_sample <= 1036263;
 925: sine_sample <= 1036508;
 926: sine_sample <= 1036750;
 927: sine_sample <= 1036990;
 928: sine_sample <= 1037227;
 929: sine_sample <= 1037462;
 930: sine_sample <= 1037694;
 931: sine_sample <= 1037924;
 932: sine_sample <= 1038151;
 933: sine_sample <= 1038376;
 934: sine_sample <= 1038599;
 935: sine_sample <= 1038819;
 936: sine_sample <= 1039037;
 937: sine_sample <= 1039252;
 938: sine_sample <= 1039465;
 939: sine_sample <= 1039675;
 940: sine_sample <= 1039883;
 941: sine_sample <= 1040089;
 942: sine_sample <= 1040292;
 943: sine_sample <= 1040492;
 944: sine_sample <= 1040690;
 945: sine_sample <= 1040886;
 946: sine_sample <= 1041079;
 947: sine_sample <= 1041270;
 948: sine_sample <= 1041458;
 949: sine_sample <= 1041644;
 950: sine_sample <= 1041828;
 951: sine_sample <= 1042009;
 952: sine_sample <= 1042187;
 953: sine_sample <= 1042363;
 954: sine_sample <= 1042537;
 955: sine_sample <= 1042708;
 956: sine_sample <= 1042877;
 957: sine_sample <= 1043043;
 958: sine_sample <= 1043207;
 959: sine_sample <= 1043368;
 960: sine_sample <= 1043527;
 961: sine_sample <= 1043683;
 962: sine_sample <= 1043837;
 963: sine_sample <= 1043989;
 964: sine_sample <= 1044138;
 965: sine_sample <= 1044285;
 966: sine_sample <= 1044429;
 967: sine_sample <= 1044570;
 968: sine_sample <= 1044710;
 969: sine_sample <= 1044846;
 970: sine_sample <= 1044981;
 971: sine_sample <= 1045113;
 972: sine_sample <= 1045242;
 973: sine_sample <= 1045369;
 974: sine_sample <= 1045493;
 975: sine_sample <= 1045615;
 976: sine_sample <= 1045735;
 977: sine_sample <= 1045852;
 978: sine_sample <= 1045967;
 979: sine_sample <= 1046079;
 980: sine_sample <= 1046189;
 981: sine_sample <= 1046296;
 982: sine_sample <= 1046401;
 983: sine_sample <= 1046503;
 984: sine_sample <= 1046603;
 985: sine_sample <= 1046700;
 986: sine_sample <= 1046795;
 987: sine_sample <= 1046888;
 988: sine_sample <= 1046978;
 989: sine_sample <= 1047065;
 990: sine_sample <= 1047150;
 991: sine_sample <= 1047233;
 992: sine_sample <= 1047313;
 993: sine_sample <= 1047391;
 994: sine_sample <= 1047466;
 995: sine_sample <= 1047539;
 996: sine_sample <= 1047609;
 997: sine_sample <= 1047677;
 998: sine_sample <= 1047742;
 999: sine_sample <= 1047805;
 1000: sine_sample <= 1047866;
 1001: sine_sample <= 1047924;
 1002: sine_sample <= 1047979;
 1003: sine_sample <= 1048032;
 1004: sine_sample <= 1048083;
 1005: sine_sample <= 1048131;
 1006: sine_sample <= 1048176;
 1007: sine_sample <= 1048220;
 1008: sine_sample <= 1048260;
 1009: sine_sample <= 1048299;
 1010: sine_sample <= 1048334;
 1011: sine_sample <= 1048368;
 1012: sine_sample <= 1048398;
 1013: sine_sample <= 1048427;
 1014: sine_sample <= 1048453;
 1015: sine_sample <= 1048476;
 1016: sine_sample <= 1048497;
 1017: sine_sample <= 1048516;
 1018: sine_sample <= 1048532;
 1019: sine_sample <= 1048545;
 1020: sine_sample <= 1048556;
 1021: sine_sample <= 1048565;
 1022: sine_sample <= 1048571;
 1023: sine_sample <= 1048575;
 1024: sine_sample <= 1048576;
 1025: sine_sample <= 1048575;
 1026: sine_sample <= 1048571;
 1027: sine_sample <= 1048565;
 1028: sine_sample <= 1048556;
 1029: sine_sample <= 1048545;
 1030: sine_sample <= 1048532;
 1031: sine_sample <= 1048516;
 1032: sine_sample <= 1048497;
 1033: sine_sample <= 1048476;
 1034: sine_sample <= 1048453;
 1035: sine_sample <= 1048427;
 1036: sine_sample <= 1048398;
 1037: sine_sample <= 1048368;
 1038: sine_sample <= 1048334;
 1039: sine_sample <= 1048299;
 1040: sine_sample <= 1048260;
 1041: sine_sample <= 1048220;
 1042: sine_sample <= 1048176;
 1043: sine_sample <= 1048131;
 1044: sine_sample <= 1048083;
 1045: sine_sample <= 1048032;
 1046: sine_sample <= 1047979;
 1047: sine_sample <= 1047924;
 1048: sine_sample <= 1047866;
 1049: sine_sample <= 1047805;
 1050: sine_sample <= 1047742;
 1051: sine_sample <= 1047677;
 1052: sine_sample <= 1047609;
 1053: sine_sample <= 1047539;
 1054: sine_sample <= 1047466;
 1055: sine_sample <= 1047391;
 1056: sine_sample <= 1047313;
 1057: sine_sample <= 1047233;
 1058: sine_sample <= 1047150;
 1059: sine_sample <= 1047065;
 1060: sine_sample <= 1046978;
 1061: sine_sample <= 1046888;
 1062: sine_sample <= 1046795;
 1063: sine_sample <= 1046700;
 1064: sine_sample <= 1046603;
 1065: sine_sample <= 1046503;
 1066: sine_sample <= 1046401;
 1067: sine_sample <= 1046296;
 1068: sine_sample <= 1046189;
 1069: sine_sample <= 1046079;
 1070: sine_sample <= 1045967;
 1071: sine_sample <= 1045852;
 1072: sine_sample <= 1045735;
 1073: sine_sample <= 1045615;
 1074: sine_sample <= 1045493;
 1075: sine_sample <= 1045369;
 1076: sine_sample <= 1045242;
 1077: sine_sample <= 1045113;
 1078: sine_sample <= 1044981;
 1079: sine_sample <= 1044846;
 1080: sine_sample <= 1044710;
 1081: sine_sample <= 1044570;
 1082: sine_sample <= 1044429;
 1083: sine_sample <= 1044285;
 1084: sine_sample <= 1044138;
 1085: sine_sample <= 1043989;
 1086: sine_sample <= 1043837;
 1087: sine_sample <= 1043683;
 1088: sine_sample <= 1043527;
 1089: sine_sample <= 1043368;
 1090: sine_sample <= 1043207;
 1091: sine_sample <= 1043043;
 1092: sine_sample <= 1042877;
 1093: sine_sample <= 1042708;
 1094: sine_sample <= 1042537;
 1095: sine_sample <= 1042363;
 1096: sine_sample <= 1042187;
 1097: sine_sample <= 1042009;
 1098: sine_sample <= 1041828;
 1099: sine_sample <= 1041644;
 1100: sine_sample <= 1041458;
 1101: sine_sample <= 1041270;
 1102: sine_sample <= 1041079;
 1103: sine_sample <= 1040886;
 1104: sine_sample <= 1040690;
 1105: sine_sample <= 1040492;
 1106: sine_sample <= 1040292;
 1107: sine_sample <= 1040089;
 1108: sine_sample <= 1039883;
 1109: sine_sample <= 1039675;
 1110: sine_sample <= 1039465;
 1111: sine_sample <= 1039252;
 1112: sine_sample <= 1039037;
 1113: sine_sample <= 1038819;
 1114: sine_sample <= 1038599;
 1115: sine_sample <= 1038376;
 1116: sine_sample <= 1038151;
 1117: sine_sample <= 1037924;
 1118: sine_sample <= 1037694;
 1119: sine_sample <= 1037462;
 1120: sine_sample <= 1037227;
 1121: sine_sample <= 1036990;
 1122: sine_sample <= 1036750;
 1123: sine_sample <= 1036508;
 1124: sine_sample <= 1036263;
 1125: sine_sample <= 1036016;
 1126: sine_sample <= 1035767;
 1127: sine_sample <= 1035515;
 1128: sine_sample <= 1035261;
 1129: sine_sample <= 1035004;
 1130: sine_sample <= 1034745;
 1131: sine_sample <= 1034483;
 1132: sine_sample <= 1034219;
 1133: sine_sample <= 1033953;
 1134: sine_sample <= 1033684;
 1135: sine_sample <= 1033412;
 1136: sine_sample <= 1033139;
 1137: sine_sample <= 1032862;
 1138: sine_sample <= 1032584;
 1139: sine_sample <= 1032303;
 1140: sine_sample <= 1032019;
 1141: sine_sample <= 1031733;
 1142: sine_sample <= 1031445;
 1143: sine_sample <= 1031154;
 1144: sine_sample <= 1030861;
 1145: sine_sample <= 1030565;
 1146: sine_sample <= 1030267;
 1147: sine_sample <= 1029967;
 1148: sine_sample <= 1029664;
 1149: sine_sample <= 1029359;
 1150: sine_sample <= 1029051;
 1151: sine_sample <= 1028741;
 1152: sine_sample <= 1028428;
 1153: sine_sample <= 1028113;
 1154: sine_sample <= 1027796;
 1155: sine_sample <= 1027476;
 1156: sine_sample <= 1027153;
 1157: sine_sample <= 1026829;
 1158: sine_sample <= 1026502;
 1159: sine_sample <= 1026172;
 1160: sine_sample <= 1025840;
 1161: sine_sample <= 1025506;
 1162: sine_sample <= 1025169;
 1163: sine_sample <= 1024830;
 1164: sine_sample <= 1024488;
 1165: sine_sample <= 1024144;
 1166: sine_sample <= 1023798;
 1167: sine_sample <= 1023449;
 1168: sine_sample <= 1023098;
 1169: sine_sample <= 1022744;
 1170: sine_sample <= 1022388;
 1171: sine_sample <= 1022030;
 1172: sine_sample <= 1021669;
 1173: sine_sample <= 1021306;
 1174: sine_sample <= 1020940;
 1175: sine_sample <= 1020572;
 1176: sine_sample <= 1020202;
 1177: sine_sample <= 1019829;
 1178: sine_sample <= 1019453;
 1179: sine_sample <= 1019076;
 1180: sine_sample <= 1018696;
 1181: sine_sample <= 1018313;
 1182: sine_sample <= 1017928;
 1183: sine_sample <= 1017541;
 1184: sine_sample <= 1017152;
 1185: sine_sample <= 1016760;
 1186: sine_sample <= 1016365;
 1187: sine_sample <= 1015968;
 1188: sine_sample <= 1015569;
 1189: sine_sample <= 1015168;
 1190: sine_sample <= 1014764;
 1191: sine_sample <= 1014357;
 1192: sine_sample <= 1013948;
 1193: sine_sample <= 1013537;
 1194: sine_sample <= 1013124;
 1195: sine_sample <= 1012708;
 1196: sine_sample <= 1012290;
 1197: sine_sample <= 1011869;
 1198: sine_sample <= 1011446;
 1199: sine_sample <= 1011020;
 1200: sine_sample <= 1010593;
 1201: sine_sample <= 1010162;
 1202: sine_sample <= 1009730;
 1203: sine_sample <= 1009295;
 1204: sine_sample <= 1008858;
 1205: sine_sample <= 1008418;
 1206: sine_sample <= 1007976;
 1207: sine_sample <= 1007531;
 1208: sine_sample <= 1007085;
 1209: sine_sample <= 1006635;
 1210: sine_sample <= 1006184;
 1211: sine_sample <= 1005730;
 1212: sine_sample <= 1005274;
 1213: sine_sample <= 1004815;
 1214: sine_sample <= 1004354;
 1215: sine_sample <= 1003891;
 1216: sine_sample <= 1003425;
 1217: sine_sample <= 1002957;
 1218: sine_sample <= 1002486;
 1219: sine_sample <= 1002013;
 1220: sine_sample <= 1001538;
 1221: sine_sample <= 1001061;
 1222: sine_sample <= 1000581;
 1223: sine_sample <= 1000099;
 1224: sine_sample <= 999614;
 1225: sine_sample <= 999127;
 1226: sine_sample <= 998638;
 1227: sine_sample <= 998146;
 1228: sine_sample <= 997652;
 1229: sine_sample <= 997156;
 1230: sine_sample <= 996657;
 1231: sine_sample <= 996156;
 1232: sine_sample <= 995653;
 1233: sine_sample <= 995147;
 1234: sine_sample <= 994639;
 1235: sine_sample <= 994128;
 1236: sine_sample <= 993616;
 1237: sine_sample <= 993101;
 1238: sine_sample <= 992583;
 1239: sine_sample <= 992063;
 1240: sine_sample <= 991541;
 1241: sine_sample <= 991017;
 1242: sine_sample <= 990490;
 1243: sine_sample <= 989961;
 1244: sine_sample <= 989430;
 1245: sine_sample <= 988896;
 1246: sine_sample <= 988360;
 1247: sine_sample <= 987821;
 1248: sine_sample <= 987281;
 1249: sine_sample <= 986738;
 1250: sine_sample <= 986192;
 1251: sine_sample <= 985645;
 1252: sine_sample <= 985095;
 1253: sine_sample <= 984542;
 1254: sine_sample <= 983988;
 1255: sine_sample <= 983431;
 1256: sine_sample <= 982871;
 1257: sine_sample <= 982310;
 1258: sine_sample <= 981746;
 1259: sine_sample <= 981180;
 1260: sine_sample <= 980611;
 1261: sine_sample <= 980040;
 1262: sine_sample <= 979467;
 1263: sine_sample <= 978892;
 1264: sine_sample <= 978314;
 1265: sine_sample <= 977734;
 1266: sine_sample <= 977152;
 1267: sine_sample <= 976567;
 1268: sine_sample <= 975980;
 1269: sine_sample <= 975391;
 1270: sine_sample <= 974799;
 1271: sine_sample <= 974205;
 1272: sine_sample <= 973609;
 1273: sine_sample <= 973011;
 1274: sine_sample <= 972410;
 1275: sine_sample <= 971807;
 1276: sine_sample <= 971202;
 1277: sine_sample <= 970594;
 1278: sine_sample <= 969985;
 1279: sine_sample <= 969372;
 1280: sine_sample <= 968758;
 1281: sine_sample <= 968141;
 1282: sine_sample <= 967522;
 1283: sine_sample <= 966901;
 1284: sine_sample <= 966278;
 1285: sine_sample <= 965652;
 1286: sine_sample <= 965024;
 1287: sine_sample <= 964393;
 1288: sine_sample <= 963761;
 1289: sine_sample <= 963126;
 1290: sine_sample <= 962489;
 1291: sine_sample <= 961849;
 1292: sine_sample <= 961208;
 1293: sine_sample <= 960564;
 1294: sine_sample <= 959918;
 1295: sine_sample <= 959269;
 1296: sine_sample <= 958619;
 1297: sine_sample <= 957966;
 1298: sine_sample <= 957310;
 1299: sine_sample <= 956653;
 1300: sine_sample <= 955993;
 1301: sine_sample <= 955331;
 1302: sine_sample <= 954667;
 1303: sine_sample <= 954001;
 1304: sine_sample <= 953332;
 1305: sine_sample <= 952661;
 1306: sine_sample <= 951988;
 1307: sine_sample <= 951312;
 1308: sine_sample <= 950635;
 1309: sine_sample <= 949955;
 1310: sine_sample <= 949273;
 1311: sine_sample <= 948588;
 1312: sine_sample <= 947902;
 1313: sine_sample <= 947213;
 1314: sine_sample <= 946522;
 1315: sine_sample <= 945828;
 1316: sine_sample <= 945133;
 1317: sine_sample <= 944435;
 1318: sine_sample <= 943735;
 1319: sine_sample <= 943033;
 1320: sine_sample <= 942329;
 1321: sine_sample <= 941622;
 1322: sine_sample <= 940913;
 1323: sine_sample <= 940202;
 1324: sine_sample <= 939489;
 1325: sine_sample <= 938773;
 1326: sine_sample <= 938056;
 1327: sine_sample <= 937336;
 1328: sine_sample <= 936614;
 1329: sine_sample <= 935889;
 1330: sine_sample <= 935163;
 1331: sine_sample <= 934434;
 1332: sine_sample <= 933703;
 1333: sine_sample <= 932970;
 1334: sine_sample <= 932235;
 1335: sine_sample <= 931497;
 1336: sine_sample <= 930758;
 1337: sine_sample <= 930016;
 1338: sine_sample <= 929272;
 1339: sine_sample <= 928526;
 1340: sine_sample <= 927777;
 1341: sine_sample <= 927027;
 1342: sine_sample <= 926274;
 1343: sine_sample <= 925519;
 1344: sine_sample <= 924762;
 1345: sine_sample <= 924002;
 1346: sine_sample <= 923241;
 1347: sine_sample <= 922477;
 1348: sine_sample <= 921711;
 1349: sine_sample <= 920943;
 1350: sine_sample <= 920173;
 1351: sine_sample <= 919401;
 1352: sine_sample <= 918626;
 1353: sine_sample <= 917850;
 1354: sine_sample <= 917071;
 1355: sine_sample <= 916290;
 1356: sine_sample <= 915507;
 1357: sine_sample <= 914721;
 1358: sine_sample <= 913934;
 1359: sine_sample <= 913144;
 1360: sine_sample <= 912352;
 1361: sine_sample <= 911559;
 1362: sine_sample <= 910763;
 1363: sine_sample <= 909964;
 1364: sine_sample <= 909164;
 1365: sine_sample <= 908362;
 1366: sine_sample <= 907557;
 1367: sine_sample <= 906750;
 1368: sine_sample <= 905941;
 1369: sine_sample <= 905130;
 1370: sine_sample <= 904317;
 1371: sine_sample <= 903502;
 1372: sine_sample <= 902685;
 1373: sine_sample <= 901865;
 1374: sine_sample <= 901043;
 1375: sine_sample <= 900220;
 1376: sine_sample <= 899394;
 1377: sine_sample <= 898566;
 1378: sine_sample <= 897736;
 1379: sine_sample <= 896903;
 1380: sine_sample <= 896069;
 1381: sine_sample <= 895233;
 1382: sine_sample <= 894394;
 1383: sine_sample <= 893553;
 1384: sine_sample <= 892711;
 1385: sine_sample <= 891866;
 1386: sine_sample <= 891019;
 1387: sine_sample <= 890170;
 1388: sine_sample <= 889319;
 1389: sine_sample <= 888466;
 1390: sine_sample <= 887610;
 1391: sine_sample <= 886753;
 1392: sine_sample <= 885893;
 1393: sine_sample <= 885032;
 1394: sine_sample <= 884168;
 1395: sine_sample <= 883302;
 1396: sine_sample <= 882434;
 1397: sine_sample <= 881565;
 1398: sine_sample <= 880693;
 1399: sine_sample <= 879819;
 1400: sine_sample <= 878942;
 1401: sine_sample <= 878064;
 1402: sine_sample <= 877184;
 1403: sine_sample <= 876302;
 1404: sine_sample <= 875417;
 1405: sine_sample <= 874531;
 1406: sine_sample <= 873642;
 1407: sine_sample <= 872752;
 1408: sine_sample <= 871859;
 1409: sine_sample <= 870965;
 1410: sine_sample <= 870068;
 1411: sine_sample <= 869169;
 1412: sine_sample <= 868268;
 1413: sine_sample <= 867365;
 1414: sine_sample <= 866461;
 1415: sine_sample <= 865554;
 1416: sine_sample <= 864645;
 1417: sine_sample <= 863734;
 1418: sine_sample <= 862821;
 1419: sine_sample <= 861906;
 1420: sine_sample <= 860989;
 1421: sine_sample <= 860069;
 1422: sine_sample <= 859148;
 1423: sine_sample <= 858225;
 1424: sine_sample <= 857300;
 1425: sine_sample <= 856373;
 1426: sine_sample <= 855444;
 1427: sine_sample <= 854512;
 1428: sine_sample <= 853579;
 1429: sine_sample <= 852644;
 1430: sine_sample <= 851707;
 1431: sine_sample <= 850767;
 1432: sine_sample <= 849826;
 1433: sine_sample <= 848883;
 1434: sine_sample <= 847938;
 1435: sine_sample <= 846990;
 1436: sine_sample <= 846041;
 1437: sine_sample <= 845090;
 1438: sine_sample <= 844137;
 1439: sine_sample <= 843181;
 1440: sine_sample <= 842224;
 1441: sine_sample <= 841265;
 1442: sine_sample <= 840304;
 1443: sine_sample <= 839341;
 1444: sine_sample <= 838376;
 1445: sine_sample <= 837409;
 1446: sine_sample <= 836440;
 1447: sine_sample <= 835469;
 1448: sine_sample <= 834496;
 1449: sine_sample <= 833521;
 1450: sine_sample <= 832544;
 1451: sine_sample <= 831565;
 1452: sine_sample <= 830584;
 1453: sine_sample <= 829601;
 1454: sine_sample <= 828617;
 1455: sine_sample <= 827630;
 1456: sine_sample <= 826641;
 1457: sine_sample <= 825651;
 1458: sine_sample <= 824658;
 1459: sine_sample <= 823664;
 1460: sine_sample <= 822667;
 1461: sine_sample <= 821669;
 1462: sine_sample <= 820669;
 1463: sine_sample <= 819667;
 1464: sine_sample <= 818662;
 1465: sine_sample <= 817656;
 1466: sine_sample <= 816648;
 1467: sine_sample <= 815639;
 1468: sine_sample <= 814627;
 1469: sine_sample <= 813613;
 1470: sine_sample <= 812597;
 1471: sine_sample <= 811580;
 1472: sine_sample <= 810560;
 1473: sine_sample <= 809539;
 1474: sine_sample <= 808516;
 1475: sine_sample <= 807491;
 1476: sine_sample <= 806463;
 1477: sine_sample <= 805434;
 1478: sine_sample <= 804404;
 1479: sine_sample <= 803371;
 1480: sine_sample <= 802336;
 1481: sine_sample <= 801300;
 1482: sine_sample <= 800261;
 1483: sine_sample <= 799221;
 1484: sine_sample <= 798179;
 1485: sine_sample <= 797135;
 1486: sine_sample <= 796089;
 1487: sine_sample <= 795041;
 1488: sine_sample <= 793991;
 1489: sine_sample <= 792940;
 1490: sine_sample <= 791886;
 1491: sine_sample <= 790831;
 1492: sine_sample <= 789774;
 1493: sine_sample <= 788715;
 1494: sine_sample <= 787654;
 1495: sine_sample <= 786591;
 1496: sine_sample <= 785527;
 1497: sine_sample <= 784460;
 1498: sine_sample <= 783392;
 1499: sine_sample <= 782322;
 1500: sine_sample <= 781250;
 1501: sine_sample <= 780176;
 1502: sine_sample <= 779100;
 1503: sine_sample <= 778023;
 1504: sine_sample <= 776944;
 1505: sine_sample <= 775863;
 1506: sine_sample <= 774780;
 1507: sine_sample <= 773695;
 1508: sine_sample <= 772608;
 1509: sine_sample <= 771520;
 1510: sine_sample <= 770430;
 1511: sine_sample <= 769338;
 1512: sine_sample <= 768244;
 1513: sine_sample <= 767148;
 1514: sine_sample <= 766051;
 1515: sine_sample <= 764951;
 1516: sine_sample <= 763850;
 1517: sine_sample <= 762748;
 1518: sine_sample <= 761643;
 1519: sine_sample <= 760536;
 1520: sine_sample <= 759428;
 1521: sine_sample <= 758318;
 1522: sine_sample <= 757206;
 1523: sine_sample <= 756093;
 1524: sine_sample <= 754977;
 1525: sine_sample <= 753860;
 1526: sine_sample <= 752741;
 1527: sine_sample <= 751621;
 1528: sine_sample <= 750498;
 1529: sine_sample <= 749374;
 1530: sine_sample <= 748248;
 1531: sine_sample <= 747120;
 1532: sine_sample <= 745991;
 1533: sine_sample <= 744860;
 1534: sine_sample <= 743727;
 1535: sine_sample <= 742592;
 1536: sine_sample <= 741455;
 1537: sine_sample <= 740317;
 1538: sine_sample <= 739177;
 1539: sine_sample <= 738035;
 1540: sine_sample <= 736892;
 1541: sine_sample <= 735747;
 1542: sine_sample <= 734600;
 1543: sine_sample <= 733451;
 1544: sine_sample <= 732301;
 1545: sine_sample <= 731149;
 1546: sine_sample <= 729995;
 1547: sine_sample <= 728839;
 1548: sine_sample <= 727682;
 1549: sine_sample <= 726523;
 1550: sine_sample <= 725362;
 1551: sine_sample <= 724200;
 1552: sine_sample <= 723036;
 1553: sine_sample <= 721870;
 1554: sine_sample <= 720702;
 1555: sine_sample <= 719533;
 1556: sine_sample <= 718362;
 1557: sine_sample <= 717190;
 1558: sine_sample <= 716016;
 1559: sine_sample <= 714840;
 1560: sine_sample <= 713662;
 1561: sine_sample <= 712483;
 1562: sine_sample <= 711302;
 1563: sine_sample <= 710119;
 1564: sine_sample <= 708935;
 1565: sine_sample <= 707749;
 1566: sine_sample <= 706561;
 1567: sine_sample <= 705372;
 1568: sine_sample <= 704181;
 1569: sine_sample <= 702988;
 1570: sine_sample <= 701794;
 1571: sine_sample <= 700598;
 1572: sine_sample <= 699400;
 1573: sine_sample <= 698201;
 1574: sine_sample <= 697000;
 1575: sine_sample <= 695798;
 1576: sine_sample <= 694593;
 1577: sine_sample <= 693388;
 1578: sine_sample <= 692180;
 1579: sine_sample <= 690971;
 1580: sine_sample <= 689760;
 1581: sine_sample <= 688548;
 1582: sine_sample <= 687334;
 1583: sine_sample <= 686119;
 1584: sine_sample <= 684901;
 1585: sine_sample <= 683683;
 1586: sine_sample <= 682462;
 1587: sine_sample <= 681240;
 1588: sine_sample <= 680017;
 1589: sine_sample <= 678792;
 1590: sine_sample <= 677565;
 1591: sine_sample <= 676336;
 1592: sine_sample <= 675106;
 1593: sine_sample <= 673875;
 1594: sine_sample <= 672642;
 1595: sine_sample <= 671407;
 1596: sine_sample <= 670171;
 1597: sine_sample <= 668933;
 1598: sine_sample <= 667693;
 1599: sine_sample <= 666452;
 1600: sine_sample <= 665210;
 1601: sine_sample <= 663966;
 1602: sine_sample <= 662720;
 1603: sine_sample <= 661473;
 1604: sine_sample <= 660224;
 1605: sine_sample <= 658973;
 1606: sine_sample <= 657721;
 1607: sine_sample <= 656468;
 1608: sine_sample <= 655213;
 1609: sine_sample <= 653956;
 1610: sine_sample <= 652698;
 1611: sine_sample <= 651438;
 1612: sine_sample <= 650177;
 1613: sine_sample <= 648915;
 1614: sine_sample <= 647650;
 1615: sine_sample <= 646384;
 1616: sine_sample <= 645117;
 1617: sine_sample <= 643848;
 1618: sine_sample <= 642578;
 1619: sine_sample <= 641306;
 1620: sine_sample <= 640033;
 1621: sine_sample <= 638758;
 1622: sine_sample <= 637482;
 1623: sine_sample <= 636204;
 1624: sine_sample <= 634924;
 1625: sine_sample <= 633644;
 1626: sine_sample <= 632361;
 1627: sine_sample <= 631077;
 1628: sine_sample <= 629792;
 1629: sine_sample <= 628505;
 1630: sine_sample <= 627217;
 1631: sine_sample <= 625927;
 1632: sine_sample <= 624636;
 1633: sine_sample <= 623343;
 1634: sine_sample <= 622049;
 1635: sine_sample <= 620754;
 1636: sine_sample <= 619457;
 1637: sine_sample <= 618158;
 1638: sine_sample <= 616858;
 1639: sine_sample <= 615557;
 1640: sine_sample <= 614254;
 1641: sine_sample <= 612949;
 1642: sine_sample <= 611644;
 1643: sine_sample <= 610336;
 1644: sine_sample <= 609028;
 1645: sine_sample <= 607718;
 1646: sine_sample <= 606406;
 1647: sine_sample <= 605093;
 1648: sine_sample <= 603779;
 1649: sine_sample <= 602463;
 1650: sine_sample <= 601146;
 1651: sine_sample <= 599827;
 1652: sine_sample <= 598507;
 1653: sine_sample <= 597186;
 1654: sine_sample <= 595863;
 1655: sine_sample <= 594539;
 1656: sine_sample <= 593213;
 1657: sine_sample <= 591886;
 1658: sine_sample <= 590557;
 1659: sine_sample <= 589228;
 1660: sine_sample <= 587896;
 1661: sine_sample <= 586564;
 1662: sine_sample <= 585230;
 1663: sine_sample <= 583894;
 1664: sine_sample <= 582558;
 1665: sine_sample <= 581220;
 1666: sine_sample <= 579880;
 1667: sine_sample <= 578539;
 1668: sine_sample <= 577197;
 1669: sine_sample <= 575854;
 1670: sine_sample <= 574509;
 1671: sine_sample <= 573162;
 1672: sine_sample <= 571815;
 1673: sine_sample <= 570466;
 1674: sine_sample <= 569116;
 1675: sine_sample <= 567764;
 1676: sine_sample <= 566411;
 1677: sine_sample <= 565057;
 1678: sine_sample <= 563701;
 1679: sine_sample <= 562344;
 1680: sine_sample <= 560986;
 1681: sine_sample <= 559626;
 1682: sine_sample <= 558265;
 1683: sine_sample <= 556903;
 1684: sine_sample <= 555539;
 1685: sine_sample <= 554175;
 1686: sine_sample <= 552808;
 1687: sine_sample <= 551441;
 1688: sine_sample <= 550072;
 1689: sine_sample <= 548702;
 1690: sine_sample <= 547331;
 1691: sine_sample <= 545958;
 1692: sine_sample <= 544584;
 1693: sine_sample <= 543209;
 1694: sine_sample <= 541833;
 1695: sine_sample <= 540455;
 1696: sine_sample <= 539076;
 1697: sine_sample <= 537696;
 1698: sine_sample <= 536314;
 1699: sine_sample <= 534931;
 1700: sine_sample <= 533547;
 1701: sine_sample <= 532162;
 1702: sine_sample <= 530775;
 1703: sine_sample <= 529387;
 1704: sine_sample <= 527998;
 1705: sine_sample <= 526608;
 1706: sine_sample <= 525217;
 1707: sine_sample <= 523824;
 1708: sine_sample <= 522430;
 1709: sine_sample <= 521034;
 1710: sine_sample <= 519638;
 1711: sine_sample <= 518240;
 1712: sine_sample <= 516841;
 1713: sine_sample <= 515441;
 1714: sine_sample <= 514040;
 1715: sine_sample <= 512637;
 1716: sine_sample <= 511234;
 1717: sine_sample <= 509829;
 1718: sine_sample <= 508422;
 1719: sine_sample <= 507015;
 1720: sine_sample <= 505606;
 1721: sine_sample <= 504197;
 1722: sine_sample <= 502786;
 1723: sine_sample <= 501374;
 1724: sine_sample <= 499960;
 1725: sine_sample <= 498546;
 1726: sine_sample <= 497130;
 1727: sine_sample <= 495713;
 1728: sine_sample <= 494295;
 1729: sine_sample <= 492876;
 1730: sine_sample <= 491456;
 1731: sine_sample <= 490035;
 1732: sine_sample <= 488612;
 1733: sine_sample <= 487188;
 1734: sine_sample <= 485763;
 1735: sine_sample <= 484337;
 1736: sine_sample <= 482910;
 1737: sine_sample <= 481482;
 1738: sine_sample <= 480052;
 1739: sine_sample <= 478622;
 1740: sine_sample <= 477190;
 1741: sine_sample <= 475757;
 1742: sine_sample <= 474323;
 1743: sine_sample <= 472888;
 1744: sine_sample <= 471452;
 1745: sine_sample <= 470014;
 1746: sine_sample <= 468576;
 1747: sine_sample <= 467137;
 1748: sine_sample <= 465696;
 1749: sine_sample <= 464254;
 1750: sine_sample <= 462811;
 1751: sine_sample <= 461368;
 1752: sine_sample <= 459923;
 1753: sine_sample <= 458477;
 1754: sine_sample <= 457029;
 1755: sine_sample <= 455581;
 1756: sine_sample <= 454132;
 1757: sine_sample <= 452682;
 1758: sine_sample <= 451230;
 1759: sine_sample <= 449778;
 1760: sine_sample <= 448324;
 1761: sine_sample <= 446870;
 1762: sine_sample <= 445414;
 1763: sine_sample <= 443957;
 1764: sine_sample <= 442499;
 1765: sine_sample <= 441041;
 1766: sine_sample <= 439581;
 1767: sine_sample <= 438120;
 1768: sine_sample <= 436658;
 1769: sine_sample <= 435195;
 1770: sine_sample <= 433731;
 1771: sine_sample <= 432266;
 1772: sine_sample <= 430800;
 1773: sine_sample <= 429333;
 1774: sine_sample <= 427865;
 1775: sine_sample <= 426396;
 1776: sine_sample <= 424926;
 1777: sine_sample <= 423455;
 1778: sine_sample <= 421983;
 1779: sine_sample <= 420510;
 1780: sine_sample <= 419036;
 1781: sine_sample <= 417562;
 1782: sine_sample <= 416086;
 1783: sine_sample <= 414609;
 1784: sine_sample <= 413131;
 1785: sine_sample <= 411652;
 1786: sine_sample <= 410172;
 1787: sine_sample <= 408691;
 1788: sine_sample <= 407209;
 1789: sine_sample <= 405727;
 1790: sine_sample <= 404243;
 1791: sine_sample <= 402758;
 1792: sine_sample <= 401273;
 1793: sine_sample <= 399786;
 1794: sine_sample <= 398299;
 1795: sine_sample <= 396810;
 1796: sine_sample <= 395321;
 1797: sine_sample <= 393831;
 1798: sine_sample <= 392340;
 1799: sine_sample <= 390847;
 1800: sine_sample <= 389354;
 1801: sine_sample <= 387860;
 1802: sine_sample <= 386366;
 1803: sine_sample <= 384870;
 1804: sine_sample <= 383373;
 1805: sine_sample <= 381876;
 1806: sine_sample <= 380377;
 1807: sine_sample <= 378878;
 1808: sine_sample <= 377377;
 1809: sine_sample <= 375876;
 1810: sine_sample <= 374374;
 1811: sine_sample <= 372871;
 1812: sine_sample <= 371367;
 1813: sine_sample <= 369863;
 1814: sine_sample <= 368357;
 1815: sine_sample <= 366851;
 1816: sine_sample <= 365344;
 1817: sine_sample <= 363835;
 1818: sine_sample <= 362326;
 1819: sine_sample <= 360817;
 1820: sine_sample <= 359306;
 1821: sine_sample <= 357794;
 1822: sine_sample <= 356282;
 1823: sine_sample <= 354769;
 1824: sine_sample <= 353255;
 1825: sine_sample <= 351740;
 1826: sine_sample <= 350224;
 1827: sine_sample <= 348708;
 1828: sine_sample <= 347190;
 1829: sine_sample <= 345672;
 1830: sine_sample <= 344153;
 1831: sine_sample <= 342633;
 1832: sine_sample <= 341113;
 1833: sine_sample <= 339591;
 1834: sine_sample <= 338069;
 1835: sine_sample <= 336546;
 1836: sine_sample <= 335022;
 1837: sine_sample <= 333498;
 1838: sine_sample <= 331972;
 1839: sine_sample <= 330446;
 1840: sine_sample <= 328919;
 1841: sine_sample <= 327392;
 1842: sine_sample <= 325863;
 1843: sine_sample <= 324334;
 1844: sine_sample <= 322804;
 1845: sine_sample <= 321273;
 1846: sine_sample <= 319742;
 1847: sine_sample <= 318209;
 1848: sine_sample <= 316676;
 1849: sine_sample <= 315143;
 1850: sine_sample <= 313608;
 1851: sine_sample <= 312073;
 1852: sine_sample <= 310537;
 1853: sine_sample <= 309000;
 1854: sine_sample <= 307463;
 1855: sine_sample <= 305925;
 1856: sine_sample <= 304386;
 1857: sine_sample <= 302846;
 1858: sine_sample <= 301306;
 1859: sine_sample <= 299765;
 1860: sine_sample <= 298223;
 1861: sine_sample <= 296681;
 1862: sine_sample <= 295138;
 1863: sine_sample <= 293594;
 1864: sine_sample <= 292049;
 1865: sine_sample <= 290504;
 1866: sine_sample <= 288958;
 1867: sine_sample <= 287412;
 1868: sine_sample <= 285864;
 1869: sine_sample <= 284316;
 1870: sine_sample <= 282768;
 1871: sine_sample <= 281219;
 1872: sine_sample <= 279669;
 1873: sine_sample <= 278118;
 1874: sine_sample <= 276567;
 1875: sine_sample <= 275015;
 1876: sine_sample <= 273463;
 1877: sine_sample <= 271909;
 1878: sine_sample <= 270356;
 1879: sine_sample <= 268801;
 1880: sine_sample <= 267246;
 1881: sine_sample <= 265690;
 1882: sine_sample <= 264134;
 1883: sine_sample <= 262577;
 1884: sine_sample <= 261020;
 1885: sine_sample <= 259461;
 1886: sine_sample <= 257903;
 1887: sine_sample <= 256343;
 1888: sine_sample <= 254783;
 1889: sine_sample <= 253223;
 1890: sine_sample <= 251662;
 1891: sine_sample <= 250100;
 1892: sine_sample <= 248537;
 1893: sine_sample <= 246974;
 1894: sine_sample <= 245411;
 1895: sine_sample <= 243847;
 1896: sine_sample <= 242282;
 1897: sine_sample <= 240717;
 1898: sine_sample <= 239151;
 1899: sine_sample <= 237585;
 1900: sine_sample <= 236018;
 1901: sine_sample <= 234450;
 1902: sine_sample <= 232882;
 1903: sine_sample <= 231314;
 1904: sine_sample <= 229744;
 1905: sine_sample <= 228175;
 1906: sine_sample <= 226605;
 1907: sine_sample <= 225034;
 1908: sine_sample <= 223462;
 1909: sine_sample <= 221891;
 1910: sine_sample <= 220318;
 1911: sine_sample <= 218746;
 1912: sine_sample <= 217172;
 1913: sine_sample <= 215598;
 1914: sine_sample <= 214024;
 1915: sine_sample <= 212449;
 1916: sine_sample <= 210874;
 1917: sine_sample <= 209298;
 1918: sine_sample <= 207721;
 1919: sine_sample <= 206145;
 1920: sine_sample <= 204567;
 1921: sine_sample <= 202989;
 1922: sine_sample <= 201411;
 1923: sine_sample <= 199832;
 1924: sine_sample <= 198253;
 1925: sine_sample <= 196673;
 1926: sine_sample <= 195093;
 1927: sine_sample <= 193512;
 1928: sine_sample <= 191931;
 1929: sine_sample <= 190350;
 1930: sine_sample <= 188768;
 1931: sine_sample <= 187185;
 1932: sine_sample <= 185603;
 1933: sine_sample <= 184019;
 1934: sine_sample <= 182435;
 1935: sine_sample <= 180851;
 1936: sine_sample <= 179267;
 1937: sine_sample <= 177682;
 1938: sine_sample <= 176096;
 1939: sine_sample <= 174510;
 1940: sine_sample <= 172924;
 1941: sine_sample <= 171337;
 1942: sine_sample <= 169750;
 1943: sine_sample <= 168163;
 1944: sine_sample <= 166575;
 1945: sine_sample <= 164987;
 1946: sine_sample <= 163398;
 1947: sine_sample <= 161809;
 1948: sine_sample <= 160220;
 1949: sine_sample <= 158630;
 1950: sine_sample <= 157040;
 1951: sine_sample <= 155449;
 1952: sine_sample <= 153858;
 1953: sine_sample <= 152267;
 1954: sine_sample <= 150675;
 1955: sine_sample <= 149083;
 1956: sine_sample <= 147491;
 1957: sine_sample <= 145898;
 1958: sine_sample <= 144305;
 1959: sine_sample <= 142712;
 1960: sine_sample <= 141118;
 1961: sine_sample <= 139524;
 1962: sine_sample <= 137930;
 1963: sine_sample <= 136335;
 1964: sine_sample <= 134740;
 1965: sine_sample <= 133145;
 1966: sine_sample <= 131549;
 1967: sine_sample <= 129953;
 1968: sine_sample <= 128357;
 1969: sine_sample <= 126760;
 1970: sine_sample <= 125164;
 1971: sine_sample <= 123566;
 1972: sine_sample <= 121969;
 1973: sine_sample <= 120371;
 1974: sine_sample <= 118773;
 1975: sine_sample <= 117175;
 1976: sine_sample <= 115576;
 1977: sine_sample <= 113978;
 1978: sine_sample <= 112379;
 1979: sine_sample <= 110779;
 1980: sine_sample <= 109180;
 1981: sine_sample <= 107580;
 1982: sine_sample <= 105980;
 1983: sine_sample <= 104379;
 1984: sine_sample <= 102779;
 1985: sine_sample <= 101178;
 1986: sine_sample <= 99577;
 1987: sine_sample <= 97975;
 1988: sine_sample <= 96374;
 1989: sine_sample <= 94772;
 1990: sine_sample <= 93170;
 1991: sine_sample <= 91568;
 1992: sine_sample <= 89965;
 1993: sine_sample <= 88362;
 1994: sine_sample <= 86760;
 1995: sine_sample <= 85156;
 1996: sine_sample <= 83553;
 1997: sine_sample <= 81950;
 1998: sine_sample <= 80346;
 1999: sine_sample <= 78742;
 2000: sine_sample <= 77138;
 2001: sine_sample <= 75534;
 2002: sine_sample <= 73930;
 2003: sine_sample <= 72325;
 2004: sine_sample <= 70720;
 2005: sine_sample <= 69115;
 2006: sine_sample <= 67510;
 2007: sine_sample <= 65905;
 2008: sine_sample <= 64300;
 2009: sine_sample <= 62694;
 2010: sine_sample <= 61088;
 2011: sine_sample <= 59483;
 2012: sine_sample <= 57877;
 2013: sine_sample <= 56270;
 2014: sine_sample <= 54664;
 2015: sine_sample <= 53058;
 2016: sine_sample <= 51451;
 2017: sine_sample <= 49845;
 2018: sine_sample <= 48238;
 2019: sine_sample <= 46631;
 2020: sine_sample <= 45024;
 2021: sine_sample <= 43417;
 2022: sine_sample <= 41810;
 2023: sine_sample <= 40203;
 2024: sine_sample <= 38595;
 2025: sine_sample <= 36988;
 2026: sine_sample <= 35380;
 2027: sine_sample <= 33773;
 2028: sine_sample <= 32165;
 2029: sine_sample <= 30557;
 2030: sine_sample <= 28949;
 2031: sine_sample <= 27341;
 2032: sine_sample <= 25733;
 2033: sine_sample <= 24125;
 2034: sine_sample <= 22517;
 2035: sine_sample <= 20909;
 2036: sine_sample <= 19301;
 2037: sine_sample <= 17693;
 2038: sine_sample <= 16084;
 2039: sine_sample <= 14476;
 2040: sine_sample <= 12868;
 2041: sine_sample <= 11259;
 2042: sine_sample <= 9651;
 2043: sine_sample <= 8043;
 2044: sine_sample <= 6434;
 2045: sine_sample <= 4826;
 2046: sine_sample <= 3217;
 2047: sine_sample <= 1609;
 2048: sine_sample <= 0;
 2049: sine_sample <= -1609;
 2050: sine_sample <= -3217;
 2051: sine_sample <= -4826;
 2052: sine_sample <= -6434;
 2053: sine_sample <= -8043;
 2054: sine_sample <= -9651;
 2055: sine_sample <= -11259;
 2056: sine_sample <= -12868;
 2057: sine_sample <= -14476;
 2058: sine_sample <= -16084;
 2059: sine_sample <= -17693;
 2060: sine_sample <= -19301;
 2061: sine_sample <= -20909;
 2062: sine_sample <= -22517;
 2063: sine_sample <= -24125;
 2064: sine_sample <= -25733;
 2065: sine_sample <= -27341;
 2066: sine_sample <= -28949;
 2067: sine_sample <= -30557;
 2068: sine_sample <= -32165;
 2069: sine_sample <= -33773;
 2070: sine_sample <= -35380;
 2071: sine_sample <= -36988;
 2072: sine_sample <= -38595;
 2073: sine_sample <= -40203;
 2074: sine_sample <= -41810;
 2075: sine_sample <= -43417;
 2076: sine_sample <= -45024;
 2077: sine_sample <= -46631;
 2078: sine_sample <= -48238;
 2079: sine_sample <= -49845;
 2080: sine_sample <= -51451;
 2081: sine_sample <= -53058;
 2082: sine_sample <= -54664;
 2083: sine_sample <= -56270;
 2084: sine_sample <= -57877;
 2085: sine_sample <= -59483;
 2086: sine_sample <= -61088;
 2087: sine_sample <= -62694;
 2088: sine_sample <= -64300;
 2089: sine_sample <= -65905;
 2090: sine_sample <= -67510;
 2091: sine_sample <= -69115;
 2092: sine_sample <= -70720;
 2093: sine_sample <= -72325;
 2094: sine_sample <= -73930;
 2095: sine_sample <= -75534;
 2096: sine_sample <= -77138;
 2097: sine_sample <= -78742;
 2098: sine_sample <= -80346;
 2099: sine_sample <= -81950;
 2100: sine_sample <= -83553;
 2101: sine_sample <= -85156;
 2102: sine_sample <= -86760;
 2103: sine_sample <= -88362;
 2104: sine_sample <= -89965;
 2105: sine_sample <= -91568;
 2106: sine_sample <= -93170;
 2107: sine_sample <= -94772;
 2108: sine_sample <= -96374;
 2109: sine_sample <= -97975;
 2110: sine_sample <= -99577;
 2111: sine_sample <= -101178;
 2112: sine_sample <= -102779;
 2113: sine_sample <= -104379;
 2114: sine_sample <= -105980;
 2115: sine_sample <= -107580;
 2116: sine_sample <= -109180;
 2117: sine_sample <= -110779;
 2118: sine_sample <= -112379;
 2119: sine_sample <= -113978;
 2120: sine_sample <= -115576;
 2121: sine_sample <= -117175;
 2122: sine_sample <= -118773;
 2123: sine_sample <= -120371;
 2124: sine_sample <= -121969;
 2125: sine_sample <= -123566;
 2126: sine_sample <= -125164;
 2127: sine_sample <= -126760;
 2128: sine_sample <= -128357;
 2129: sine_sample <= -129953;
 2130: sine_sample <= -131549;
 2131: sine_sample <= -133145;
 2132: sine_sample <= -134740;
 2133: sine_sample <= -136335;
 2134: sine_sample <= -137930;
 2135: sine_sample <= -139524;
 2136: sine_sample <= -141118;
 2137: sine_sample <= -142712;
 2138: sine_sample <= -144305;
 2139: sine_sample <= -145898;
 2140: sine_sample <= -147491;
 2141: sine_sample <= -149083;
 2142: sine_sample <= -150675;
 2143: sine_sample <= -152267;
 2144: sine_sample <= -153858;
 2145: sine_sample <= -155449;
 2146: sine_sample <= -157040;
 2147: sine_sample <= -158630;
 2148: sine_sample <= -160220;
 2149: sine_sample <= -161809;
 2150: sine_sample <= -163398;
 2151: sine_sample <= -164987;
 2152: sine_sample <= -166575;
 2153: sine_sample <= -168163;
 2154: sine_sample <= -169750;
 2155: sine_sample <= -171337;
 2156: sine_sample <= -172924;
 2157: sine_sample <= -174510;
 2158: sine_sample <= -176096;
 2159: sine_sample <= -177682;
 2160: sine_sample <= -179267;
 2161: sine_sample <= -180851;
 2162: sine_sample <= -182435;
 2163: sine_sample <= -184019;
 2164: sine_sample <= -185603;
 2165: sine_sample <= -187185;
 2166: sine_sample <= -188768;
 2167: sine_sample <= -190350;
 2168: sine_sample <= -191931;
 2169: sine_sample <= -193512;
 2170: sine_sample <= -195093;
 2171: sine_sample <= -196673;
 2172: sine_sample <= -198253;
 2173: sine_sample <= -199832;
 2174: sine_sample <= -201411;
 2175: sine_sample <= -202989;
 2176: sine_sample <= -204567;
 2177: sine_sample <= -206145;
 2178: sine_sample <= -207721;
 2179: sine_sample <= -209298;
 2180: sine_sample <= -210874;
 2181: sine_sample <= -212449;
 2182: sine_sample <= -214024;
 2183: sine_sample <= -215598;
 2184: sine_sample <= -217172;
 2185: sine_sample <= -218746;
 2186: sine_sample <= -220318;
 2187: sine_sample <= -221891;
 2188: sine_sample <= -223462;
 2189: sine_sample <= -225034;
 2190: sine_sample <= -226605;
 2191: sine_sample <= -228175;
 2192: sine_sample <= -229744;
 2193: sine_sample <= -231314;
 2194: sine_sample <= -232882;
 2195: sine_sample <= -234450;
 2196: sine_sample <= -236018;
 2197: sine_sample <= -237585;
 2198: sine_sample <= -239151;
 2199: sine_sample <= -240717;
 2200: sine_sample <= -242282;
 2201: sine_sample <= -243847;
 2202: sine_sample <= -245411;
 2203: sine_sample <= -246974;
 2204: sine_sample <= -248537;
 2205: sine_sample <= -250100;
 2206: sine_sample <= -251662;
 2207: sine_sample <= -253223;
 2208: sine_sample <= -254783;
 2209: sine_sample <= -256343;
 2210: sine_sample <= -257903;
 2211: sine_sample <= -259461;
 2212: sine_sample <= -261020;
 2213: sine_sample <= -262577;
 2214: sine_sample <= -264134;
 2215: sine_sample <= -265690;
 2216: sine_sample <= -267246;
 2217: sine_sample <= -268801;
 2218: sine_sample <= -270356;
 2219: sine_sample <= -271909;
 2220: sine_sample <= -273463;
 2221: sine_sample <= -275015;
 2222: sine_sample <= -276567;
 2223: sine_sample <= -278118;
 2224: sine_sample <= -279669;
 2225: sine_sample <= -281219;
 2226: sine_sample <= -282768;
 2227: sine_sample <= -284316;
 2228: sine_sample <= -285864;
 2229: sine_sample <= -287412;
 2230: sine_sample <= -288958;
 2231: sine_sample <= -290504;
 2232: sine_sample <= -292049;
 2233: sine_sample <= -293594;
 2234: sine_sample <= -295138;
 2235: sine_sample <= -296681;
 2236: sine_sample <= -298223;
 2237: sine_sample <= -299765;
 2238: sine_sample <= -301306;
 2239: sine_sample <= -302846;
 2240: sine_sample <= -304386;
 2241: sine_sample <= -305925;
 2242: sine_sample <= -307463;
 2243: sine_sample <= -309000;
 2244: sine_sample <= -310537;
 2245: sine_sample <= -312073;
 2246: sine_sample <= -313608;
 2247: sine_sample <= -315143;
 2248: sine_sample <= -316676;
 2249: sine_sample <= -318209;
 2250: sine_sample <= -319742;
 2251: sine_sample <= -321273;
 2252: sine_sample <= -322804;
 2253: sine_sample <= -324334;
 2254: sine_sample <= -325863;
 2255: sine_sample <= -327392;
 2256: sine_sample <= -328919;
 2257: sine_sample <= -330446;
 2258: sine_sample <= -331972;
 2259: sine_sample <= -333498;
 2260: sine_sample <= -335022;
 2261: sine_sample <= -336546;
 2262: sine_sample <= -338069;
 2263: sine_sample <= -339591;
 2264: sine_sample <= -341113;
 2265: sine_sample <= -342633;
 2266: sine_sample <= -344153;
 2267: sine_sample <= -345672;
 2268: sine_sample <= -347190;
 2269: sine_sample <= -348708;
 2270: sine_sample <= -350224;
 2271: sine_sample <= -351740;
 2272: sine_sample <= -353255;
 2273: sine_sample <= -354769;
 2274: sine_sample <= -356282;
 2275: sine_sample <= -357794;
 2276: sine_sample <= -359306;
 2277: sine_sample <= -360817;
 2278: sine_sample <= -362326;
 2279: sine_sample <= -363835;
 2280: sine_sample <= -365344;
 2281: sine_sample <= -366851;
 2282: sine_sample <= -368357;
 2283: sine_sample <= -369863;
 2284: sine_sample <= -371367;
 2285: sine_sample <= -372871;
 2286: sine_sample <= -374374;
 2287: sine_sample <= -375876;
 2288: sine_sample <= -377377;
 2289: sine_sample <= -378878;
 2290: sine_sample <= -380377;
 2291: sine_sample <= -381876;
 2292: sine_sample <= -383373;
 2293: sine_sample <= -384870;
 2294: sine_sample <= -386366;
 2295: sine_sample <= -387860;
 2296: sine_sample <= -389354;
 2297: sine_sample <= -390847;
 2298: sine_sample <= -392340;
 2299: sine_sample <= -393831;
 2300: sine_sample <= -395321;
 2301: sine_sample <= -396810;
 2302: sine_sample <= -398299;
 2303: sine_sample <= -399786;
 2304: sine_sample <= -401273;
 2305: sine_sample <= -402758;
 2306: sine_sample <= -404243;
 2307: sine_sample <= -405727;
 2308: sine_sample <= -407209;
 2309: sine_sample <= -408691;
 2310: sine_sample <= -410172;
 2311: sine_sample <= -411652;
 2312: sine_sample <= -413131;
 2313: sine_sample <= -414609;
 2314: sine_sample <= -416086;
 2315: sine_sample <= -417562;
 2316: sine_sample <= -419036;
 2317: sine_sample <= -420510;
 2318: sine_sample <= -421983;
 2319: sine_sample <= -423455;
 2320: sine_sample <= -424926;
 2321: sine_sample <= -426396;
 2322: sine_sample <= -427865;
 2323: sine_sample <= -429333;
 2324: sine_sample <= -430800;
 2325: sine_sample <= -432266;
 2326: sine_sample <= -433731;
 2327: sine_sample <= -435195;
 2328: sine_sample <= -436658;
 2329: sine_sample <= -438120;
 2330: sine_sample <= -439581;
 2331: sine_sample <= -441041;
 2332: sine_sample <= -442499;
 2333: sine_sample <= -443957;
 2334: sine_sample <= -445414;
 2335: sine_sample <= -446870;
 2336: sine_sample <= -448324;
 2337: sine_sample <= -449778;
 2338: sine_sample <= -451230;
 2339: sine_sample <= -452682;
 2340: sine_sample <= -454132;
 2341: sine_sample <= -455581;
 2342: sine_sample <= -457029;
 2343: sine_sample <= -458477;
 2344: sine_sample <= -459923;
 2345: sine_sample <= -461368;
 2346: sine_sample <= -462811;
 2347: sine_sample <= -464254;
 2348: sine_sample <= -465696;
 2349: sine_sample <= -467137;
 2350: sine_sample <= -468576;
 2351: sine_sample <= -470014;
 2352: sine_sample <= -471452;
 2353: sine_sample <= -472888;
 2354: sine_sample <= -474323;
 2355: sine_sample <= -475757;
 2356: sine_sample <= -477190;
 2357: sine_sample <= -478622;
 2358: sine_sample <= -480052;
 2359: sine_sample <= -481482;
 2360: sine_sample <= -482910;
 2361: sine_sample <= -484337;
 2362: sine_sample <= -485763;
 2363: sine_sample <= -487188;
 2364: sine_sample <= -488612;
 2365: sine_sample <= -490035;
 2366: sine_sample <= -491456;
 2367: sine_sample <= -492876;
 2368: sine_sample <= -494295;
 2369: sine_sample <= -495713;
 2370: sine_sample <= -497130;
 2371: sine_sample <= -498546;
 2372: sine_sample <= -499960;
 2373: sine_sample <= -501374;
 2374: sine_sample <= -502786;
 2375: sine_sample <= -504197;
 2376: sine_sample <= -505606;
 2377: sine_sample <= -507015;
 2378: sine_sample <= -508422;
 2379: sine_sample <= -509829;
 2380: sine_sample <= -511234;
 2381: sine_sample <= -512637;
 2382: sine_sample <= -514040;
 2383: sine_sample <= -515441;
 2384: sine_sample <= -516841;
 2385: sine_sample <= -518240;
 2386: sine_sample <= -519638;
 2387: sine_sample <= -521034;
 2388: sine_sample <= -522430;
 2389: sine_sample <= -523824;
 2390: sine_sample <= -525217;
 2391: sine_sample <= -526608;
 2392: sine_sample <= -527998;
 2393: sine_sample <= -529387;
 2394: sine_sample <= -530775;
 2395: sine_sample <= -532162;
 2396: sine_sample <= -533547;
 2397: sine_sample <= -534931;
 2398: sine_sample <= -536314;
 2399: sine_sample <= -537696;
 2400: sine_sample <= -539076;
 2401: sine_sample <= -540455;
 2402: sine_sample <= -541833;
 2403: sine_sample <= -543209;
 2404: sine_sample <= -544584;
 2405: sine_sample <= -545958;
 2406: sine_sample <= -547331;
 2407: sine_sample <= -548702;
 2408: sine_sample <= -550072;
 2409: sine_sample <= -551441;
 2410: sine_sample <= -552808;
 2411: sine_sample <= -554175;
 2412: sine_sample <= -555539;
 2413: sine_sample <= -556903;
 2414: sine_sample <= -558265;
 2415: sine_sample <= -559626;
 2416: sine_sample <= -560986;
 2417: sine_sample <= -562344;
 2418: sine_sample <= -563701;
 2419: sine_sample <= -565057;
 2420: sine_sample <= -566411;
 2421: sine_sample <= -567764;
 2422: sine_sample <= -569116;
 2423: sine_sample <= -570466;
 2424: sine_sample <= -571815;
 2425: sine_sample <= -573162;
 2426: sine_sample <= -574509;
 2427: sine_sample <= -575854;
 2428: sine_sample <= -577197;
 2429: sine_sample <= -578539;
 2430: sine_sample <= -579880;
 2431: sine_sample <= -581220;
 2432: sine_sample <= -582558;
 2433: sine_sample <= -583894;
 2434: sine_sample <= -585230;
 2435: sine_sample <= -586564;
 2436: sine_sample <= -587896;
 2437: sine_sample <= -589228;
 2438: sine_sample <= -590557;
 2439: sine_sample <= -591886;
 2440: sine_sample <= -593213;
 2441: sine_sample <= -594539;
 2442: sine_sample <= -595863;
 2443: sine_sample <= -597186;
 2444: sine_sample <= -598507;
 2445: sine_sample <= -599827;
 2446: sine_sample <= -601146;
 2447: sine_sample <= -602463;
 2448: sine_sample <= -603779;
 2449: sine_sample <= -605093;
 2450: sine_sample <= -606406;
 2451: sine_sample <= -607718;
 2452: sine_sample <= -609028;
 2453: sine_sample <= -610336;
 2454: sine_sample <= -611644;
 2455: sine_sample <= -612949;
 2456: sine_sample <= -614254;
 2457: sine_sample <= -615557;
 2458: sine_sample <= -616858;
 2459: sine_sample <= -618158;
 2460: sine_sample <= -619457;
 2461: sine_sample <= -620754;
 2462: sine_sample <= -622049;
 2463: sine_sample <= -623343;
 2464: sine_sample <= -624636;
 2465: sine_sample <= -625927;
 2466: sine_sample <= -627217;
 2467: sine_sample <= -628505;
 2468: sine_sample <= -629792;
 2469: sine_sample <= -631077;
 2470: sine_sample <= -632361;
 2471: sine_sample <= -633644;
 2472: sine_sample <= -634924;
 2473: sine_sample <= -636204;
 2474: sine_sample <= -637482;
 2475: sine_sample <= -638758;
 2476: sine_sample <= -640033;
 2477: sine_sample <= -641306;
 2478: sine_sample <= -642578;
 2479: sine_sample <= -643848;
 2480: sine_sample <= -645117;
 2481: sine_sample <= -646384;
 2482: sine_sample <= -647650;
 2483: sine_sample <= -648915;
 2484: sine_sample <= -650177;
 2485: sine_sample <= -651438;
 2486: sine_sample <= -652698;
 2487: sine_sample <= -653956;
 2488: sine_sample <= -655213;
 2489: sine_sample <= -656468;
 2490: sine_sample <= -657721;
 2491: sine_sample <= -658973;
 2492: sine_sample <= -660224;
 2493: sine_sample <= -661473;
 2494: sine_sample <= -662720;
 2495: sine_sample <= -663966;
 2496: sine_sample <= -665210;
 2497: sine_sample <= -666452;
 2498: sine_sample <= -667693;
 2499: sine_sample <= -668933;
 2500: sine_sample <= -670171;
 2501: sine_sample <= -671407;
 2502: sine_sample <= -672642;
 2503: sine_sample <= -673875;
 2504: sine_sample <= -675106;
 2505: sine_sample <= -676336;
 2506: sine_sample <= -677565;
 2507: sine_sample <= -678792;
 2508: sine_sample <= -680017;
 2509: sine_sample <= -681240;
 2510: sine_sample <= -682462;
 2511: sine_sample <= -683683;
 2512: sine_sample <= -684901;
 2513: sine_sample <= -686119;
 2514: sine_sample <= -687334;
 2515: sine_sample <= -688548;
 2516: sine_sample <= -689760;
 2517: sine_sample <= -690971;
 2518: sine_sample <= -692180;
 2519: sine_sample <= -693388;
 2520: sine_sample <= -694593;
 2521: sine_sample <= -695798;
 2522: sine_sample <= -697000;
 2523: sine_sample <= -698201;
 2524: sine_sample <= -699400;
 2525: sine_sample <= -700598;
 2526: sine_sample <= -701794;
 2527: sine_sample <= -702988;
 2528: sine_sample <= -704181;
 2529: sine_sample <= -705372;
 2530: sine_sample <= -706561;
 2531: sine_sample <= -707749;
 2532: sine_sample <= -708935;
 2533: sine_sample <= -710119;
 2534: sine_sample <= -711302;
 2535: sine_sample <= -712483;
 2536: sine_sample <= -713662;
 2537: sine_sample <= -714840;
 2538: sine_sample <= -716016;
 2539: sine_sample <= -717190;
 2540: sine_sample <= -718362;
 2541: sine_sample <= -719533;
 2542: sine_sample <= -720702;
 2543: sine_sample <= -721870;
 2544: sine_sample <= -723036;
 2545: sine_sample <= -724200;
 2546: sine_sample <= -725362;
 2547: sine_sample <= -726523;
 2548: sine_sample <= -727682;
 2549: sine_sample <= -728839;
 2550: sine_sample <= -729995;
 2551: sine_sample <= -731149;
 2552: sine_sample <= -732301;
 2553: sine_sample <= -733451;
 2554: sine_sample <= -734600;
 2555: sine_sample <= -735747;
 2556: sine_sample <= -736892;
 2557: sine_sample <= -738035;
 2558: sine_sample <= -739177;
 2559: sine_sample <= -740317;
 2560: sine_sample <= -741455;
 2561: sine_sample <= -742592;
 2562: sine_sample <= -743727;
 2563: sine_sample <= -744860;
 2564: sine_sample <= -745991;
 2565: sine_sample <= -747120;
 2566: sine_sample <= -748248;
 2567: sine_sample <= -749374;
 2568: sine_sample <= -750498;
 2569: sine_sample <= -751621;
 2570: sine_sample <= -752741;
 2571: sine_sample <= -753860;
 2572: sine_sample <= -754977;
 2573: sine_sample <= -756093;
 2574: sine_sample <= -757206;
 2575: sine_sample <= -758318;
 2576: sine_sample <= -759428;
 2577: sine_sample <= -760536;
 2578: sine_sample <= -761643;
 2579: sine_sample <= -762748;
 2580: sine_sample <= -763850;
 2581: sine_sample <= -764951;
 2582: sine_sample <= -766051;
 2583: sine_sample <= -767148;
 2584: sine_sample <= -768244;
 2585: sine_sample <= -769338;
 2586: sine_sample <= -770430;
 2587: sine_sample <= -771520;
 2588: sine_sample <= -772608;
 2589: sine_sample <= -773695;
 2590: sine_sample <= -774780;
 2591: sine_sample <= -775863;
 2592: sine_sample <= -776944;
 2593: sine_sample <= -778023;
 2594: sine_sample <= -779100;
 2595: sine_sample <= -780176;
 2596: sine_sample <= -781250;
 2597: sine_sample <= -782322;
 2598: sine_sample <= -783392;
 2599: sine_sample <= -784460;
 2600: sine_sample <= -785527;
 2601: sine_sample <= -786591;
 2602: sine_sample <= -787654;
 2603: sine_sample <= -788715;
 2604: sine_sample <= -789774;
 2605: sine_sample <= -790831;
 2606: sine_sample <= -791886;
 2607: sine_sample <= -792940;
 2608: sine_sample <= -793991;
 2609: sine_sample <= -795041;
 2610: sine_sample <= -796089;
 2611: sine_sample <= -797135;
 2612: sine_sample <= -798179;
 2613: sine_sample <= -799221;
 2614: sine_sample <= -800261;
 2615: sine_sample <= -801300;
 2616: sine_sample <= -802336;
 2617: sine_sample <= -803371;
 2618: sine_sample <= -804404;
 2619: sine_sample <= -805434;
 2620: sine_sample <= -806463;
 2621: sine_sample <= -807491;
 2622: sine_sample <= -808516;
 2623: sine_sample <= -809539;
 2624: sine_sample <= -810560;
 2625: sine_sample <= -811580;
 2626: sine_sample <= -812597;
 2627: sine_sample <= -813613;
 2628: sine_sample <= -814627;
 2629: sine_sample <= -815639;
 2630: sine_sample <= -816648;
 2631: sine_sample <= -817656;
 2632: sine_sample <= -818662;
 2633: sine_sample <= -819667;
 2634: sine_sample <= -820669;
 2635: sine_sample <= -821669;
 2636: sine_sample <= -822667;
 2637: sine_sample <= -823664;
 2638: sine_sample <= -824658;
 2639: sine_sample <= -825651;
 2640: sine_sample <= -826641;
 2641: sine_sample <= -827630;
 2642: sine_sample <= -828617;
 2643: sine_sample <= -829601;
 2644: sine_sample <= -830584;
 2645: sine_sample <= -831565;
 2646: sine_sample <= -832544;
 2647: sine_sample <= -833521;
 2648: sine_sample <= -834496;
 2649: sine_sample <= -835469;
 2650: sine_sample <= -836440;
 2651: sine_sample <= -837409;
 2652: sine_sample <= -838376;
 2653: sine_sample <= -839341;
 2654: sine_sample <= -840304;
 2655: sine_sample <= -841265;
 2656: sine_sample <= -842224;
 2657: sine_sample <= -843181;
 2658: sine_sample <= -844137;
 2659: sine_sample <= -845090;
 2660: sine_sample <= -846041;
 2661: sine_sample <= -846990;
 2662: sine_sample <= -847938;
 2663: sine_sample <= -848883;
 2664: sine_sample <= -849826;
 2665: sine_sample <= -850767;
 2666: sine_sample <= -851707;
 2667: sine_sample <= -852644;
 2668: sine_sample <= -853579;
 2669: sine_sample <= -854512;
 2670: sine_sample <= -855444;
 2671: sine_sample <= -856373;
 2672: sine_sample <= -857300;
 2673: sine_sample <= -858225;
 2674: sine_sample <= -859148;
 2675: sine_sample <= -860069;
 2676: sine_sample <= -860989;
 2677: sine_sample <= -861906;
 2678: sine_sample <= -862821;
 2679: sine_sample <= -863734;
 2680: sine_sample <= -864645;
 2681: sine_sample <= -865554;
 2682: sine_sample <= -866461;
 2683: sine_sample <= -867365;
 2684: sine_sample <= -868268;
 2685: sine_sample <= -869169;
 2686: sine_sample <= -870068;
 2687: sine_sample <= -870965;
 2688: sine_sample <= -871859;
 2689: sine_sample <= -872752;
 2690: sine_sample <= -873642;
 2691: sine_sample <= -874531;
 2692: sine_sample <= -875417;
 2693: sine_sample <= -876302;
 2694: sine_sample <= -877184;
 2695: sine_sample <= -878064;
 2696: sine_sample <= -878942;
 2697: sine_sample <= -879819;
 2698: sine_sample <= -880693;
 2699: sine_sample <= -881565;
 2700: sine_sample <= -882434;
 2701: sine_sample <= -883302;
 2702: sine_sample <= -884168;
 2703: sine_sample <= -885032;
 2704: sine_sample <= -885893;
 2705: sine_sample <= -886753;
 2706: sine_sample <= -887610;
 2707: sine_sample <= -888466;
 2708: sine_sample <= -889319;
 2709: sine_sample <= -890170;
 2710: sine_sample <= -891019;
 2711: sine_sample <= -891866;
 2712: sine_sample <= -892711;
 2713: sine_sample <= -893553;
 2714: sine_sample <= -894394;
 2715: sine_sample <= -895233;
 2716: sine_sample <= -896069;
 2717: sine_sample <= -896903;
 2718: sine_sample <= -897736;
 2719: sine_sample <= -898566;
 2720: sine_sample <= -899394;
 2721: sine_sample <= -900220;
 2722: sine_sample <= -901043;
 2723: sine_sample <= -901865;
 2724: sine_sample <= -902685;
 2725: sine_sample <= -903502;
 2726: sine_sample <= -904317;
 2727: sine_sample <= -905130;
 2728: sine_sample <= -905941;
 2729: sine_sample <= -906750;
 2730: sine_sample <= -907557;
 2731: sine_sample <= -908362;
 2732: sine_sample <= -909164;
 2733: sine_sample <= -909964;
 2734: sine_sample <= -910763;
 2735: sine_sample <= -911559;
 2736: sine_sample <= -912352;
 2737: sine_sample <= -913144;
 2738: sine_sample <= -913934;
 2739: sine_sample <= -914721;
 2740: sine_sample <= -915507;
 2741: sine_sample <= -916290;
 2742: sine_sample <= -917071;
 2743: sine_sample <= -917850;
 2744: sine_sample <= -918626;
 2745: sine_sample <= -919401;
 2746: sine_sample <= -920173;
 2747: sine_sample <= -920943;
 2748: sine_sample <= -921711;
 2749: sine_sample <= -922477;
 2750: sine_sample <= -923241;
 2751: sine_sample <= -924002;
 2752: sine_sample <= -924762;
 2753: sine_sample <= -925519;
 2754: sine_sample <= -926274;
 2755: sine_sample <= -927027;
 2756: sine_sample <= -927777;
 2757: sine_sample <= -928526;
 2758: sine_sample <= -929272;
 2759: sine_sample <= -930016;
 2760: sine_sample <= -930758;
 2761: sine_sample <= -931497;
 2762: sine_sample <= -932235;
 2763: sine_sample <= -932970;
 2764: sine_sample <= -933703;
 2765: sine_sample <= -934434;
 2766: sine_sample <= -935163;
 2767: sine_sample <= -935889;
 2768: sine_sample <= -936614;
 2769: sine_sample <= -937336;
 2770: sine_sample <= -938056;
 2771: sine_sample <= -938773;
 2772: sine_sample <= -939489;
 2773: sine_sample <= -940202;
 2774: sine_sample <= -940913;
 2775: sine_sample <= -941622;
 2776: sine_sample <= -942329;
 2777: sine_sample <= -943033;
 2778: sine_sample <= -943735;
 2779: sine_sample <= -944435;
 2780: sine_sample <= -945133;
 2781: sine_sample <= -945828;
 2782: sine_sample <= -946522;
 2783: sine_sample <= -947213;
 2784: sine_sample <= -947902;
 2785: sine_sample <= -948588;
 2786: sine_sample <= -949273;
 2787: sine_sample <= -949955;
 2788: sine_sample <= -950635;
 2789: sine_sample <= -951312;
 2790: sine_sample <= -951988;
 2791: sine_sample <= -952661;
 2792: sine_sample <= -953332;
 2793: sine_sample <= -954001;
 2794: sine_sample <= -954667;
 2795: sine_sample <= -955331;
 2796: sine_sample <= -955993;
 2797: sine_sample <= -956653;
 2798: sine_sample <= -957310;
 2799: sine_sample <= -957966;
 2800: sine_sample <= -958619;
 2801: sine_sample <= -959269;
 2802: sine_sample <= -959918;
 2803: sine_sample <= -960564;
 2804: sine_sample <= -961208;
 2805: sine_sample <= -961849;
 2806: sine_sample <= -962489;
 2807: sine_sample <= -963126;
 2808: sine_sample <= -963761;
 2809: sine_sample <= -964393;
 2810: sine_sample <= -965024;
 2811: sine_sample <= -965652;
 2812: sine_sample <= -966278;
 2813: sine_sample <= -966901;
 2814: sine_sample <= -967522;
 2815: sine_sample <= -968141;
 2816: sine_sample <= -968758;
 2817: sine_sample <= -969372;
 2818: sine_sample <= -969985;
 2819: sine_sample <= -970594;
 2820: sine_sample <= -971202;
 2821: sine_sample <= -971807;
 2822: sine_sample <= -972410;
 2823: sine_sample <= -973011;
 2824: sine_sample <= -973609;
 2825: sine_sample <= -974205;
 2826: sine_sample <= -974799;
 2827: sine_sample <= -975391;
 2828: sine_sample <= -975980;
 2829: sine_sample <= -976567;
 2830: sine_sample <= -977152;
 2831: sine_sample <= -977734;
 2832: sine_sample <= -978314;
 2833: sine_sample <= -978892;
 2834: sine_sample <= -979467;
 2835: sine_sample <= -980040;
 2836: sine_sample <= -980611;
 2837: sine_sample <= -981180;
 2838: sine_sample <= -981746;
 2839: sine_sample <= -982310;
 2840: sine_sample <= -982871;
 2841: sine_sample <= -983431;
 2842: sine_sample <= -983988;
 2843: sine_sample <= -984542;
 2844: sine_sample <= -985095;
 2845: sine_sample <= -985645;
 2846: sine_sample <= -986192;
 2847: sine_sample <= -986738;
 2848: sine_sample <= -987281;
 2849: sine_sample <= -987821;
 2850: sine_sample <= -988360;
 2851: sine_sample <= -988896;
 2852: sine_sample <= -989430;
 2853: sine_sample <= -989961;
 2854: sine_sample <= -990490;
 2855: sine_sample <= -991017;
 2856: sine_sample <= -991541;
 2857: sine_sample <= -992063;
 2858: sine_sample <= -992583;
 2859: sine_sample <= -993101;
 2860: sine_sample <= -993616;
 2861: sine_sample <= -994128;
 2862: sine_sample <= -994639;
 2863: sine_sample <= -995147;
 2864: sine_sample <= -995653;
 2865: sine_sample <= -996156;
 2866: sine_sample <= -996657;
 2867: sine_sample <= -997156;
 2868: sine_sample <= -997652;
 2869: sine_sample <= -998146;
 2870: sine_sample <= -998638;
 2871: sine_sample <= -999127;
 2872: sine_sample <= -999614;
 2873: sine_sample <= -1000099;
 2874: sine_sample <= -1000581;
 2875: sine_sample <= -1001061;
 2876: sine_sample <= -1001538;
 2877: sine_sample <= -1002013;
 2878: sine_sample <= -1002486;
 2879: sine_sample <= -1002957;
 2880: sine_sample <= -1003425;
 2881: sine_sample <= -1003891;
 2882: sine_sample <= -1004354;
 2883: sine_sample <= -1004815;
 2884: sine_sample <= -1005274;
 2885: sine_sample <= -1005730;
 2886: sine_sample <= -1006184;
 2887: sine_sample <= -1006635;
 2888: sine_sample <= -1007085;
 2889: sine_sample <= -1007531;
 2890: sine_sample <= -1007976;
 2891: sine_sample <= -1008418;
 2892: sine_sample <= -1008858;
 2893: sine_sample <= -1009295;
 2894: sine_sample <= -1009730;
 2895: sine_sample <= -1010162;
 2896: sine_sample <= -1010593;
 2897: sine_sample <= -1011020;
 2898: sine_sample <= -1011446;
 2899: sine_sample <= -1011869;
 2900: sine_sample <= -1012290;
 2901: sine_sample <= -1012708;
 2902: sine_sample <= -1013124;
 2903: sine_sample <= -1013537;
 2904: sine_sample <= -1013948;
 2905: sine_sample <= -1014357;
 2906: sine_sample <= -1014764;
 2907: sine_sample <= -1015168;
 2908: sine_sample <= -1015569;
 2909: sine_sample <= -1015968;
 2910: sine_sample <= -1016365;
 2911: sine_sample <= -1016760;
 2912: sine_sample <= -1017152;
 2913: sine_sample <= -1017541;
 2914: sine_sample <= -1017928;
 2915: sine_sample <= -1018313;
 2916: sine_sample <= -1018696;
 2917: sine_sample <= -1019076;
 2918: sine_sample <= -1019453;
 2919: sine_sample <= -1019829;
 2920: sine_sample <= -1020202;
 2921: sine_sample <= -1020572;
 2922: sine_sample <= -1020940;
 2923: sine_sample <= -1021306;
 2924: sine_sample <= -1021669;
 2925: sine_sample <= -1022030;
 2926: sine_sample <= -1022388;
 2927: sine_sample <= -1022744;
 2928: sine_sample <= -1023098;
 2929: sine_sample <= -1023449;
 2930: sine_sample <= -1023798;
 2931: sine_sample <= -1024144;
 2932: sine_sample <= -1024488;
 2933: sine_sample <= -1024830;
 2934: sine_sample <= -1025169;
 2935: sine_sample <= -1025506;
 2936: sine_sample <= -1025840;
 2937: sine_sample <= -1026172;
 2938: sine_sample <= -1026502;
 2939: sine_sample <= -1026829;
 2940: sine_sample <= -1027153;
 2941: sine_sample <= -1027476;
 2942: sine_sample <= -1027796;
 2943: sine_sample <= -1028113;
 2944: sine_sample <= -1028428;
 2945: sine_sample <= -1028741;
 2946: sine_sample <= -1029051;
 2947: sine_sample <= -1029359;
 2948: sine_sample <= -1029664;
 2949: sine_sample <= -1029967;
 2950: sine_sample <= -1030267;
 2951: sine_sample <= -1030565;
 2952: sine_sample <= -1030861;
 2953: sine_sample <= -1031154;
 2954: sine_sample <= -1031445;
 2955: sine_sample <= -1031733;
 2956: sine_sample <= -1032019;
 2957: sine_sample <= -1032303;
 2958: sine_sample <= -1032584;
 2959: sine_sample <= -1032862;
 2960: sine_sample <= -1033139;
 2961: sine_sample <= -1033412;
 2962: sine_sample <= -1033684;
 2963: sine_sample <= -1033953;
 2964: sine_sample <= -1034219;
 2965: sine_sample <= -1034483;
 2966: sine_sample <= -1034745;
 2967: sine_sample <= -1035004;
 2968: sine_sample <= -1035261;
 2969: sine_sample <= -1035515;
 2970: sine_sample <= -1035767;
 2971: sine_sample <= -1036016;
 2972: sine_sample <= -1036263;
 2973: sine_sample <= -1036508;
 2974: sine_sample <= -1036750;
 2975: sine_sample <= -1036990;
 2976: sine_sample <= -1037227;
 2977: sine_sample <= -1037462;
 2978: sine_sample <= -1037694;
 2979: sine_sample <= -1037924;
 2980: sine_sample <= -1038151;
 2981: sine_sample <= -1038376;
 2982: sine_sample <= -1038599;
 2983: sine_sample <= -1038819;
 2984: sine_sample <= -1039037;
 2985: sine_sample <= -1039252;
 2986: sine_sample <= -1039465;
 2987: sine_sample <= -1039675;
 2988: sine_sample <= -1039883;
 2989: sine_sample <= -1040089;
 2990: sine_sample <= -1040292;
 2991: sine_sample <= -1040492;
 2992: sine_sample <= -1040690;
 2993: sine_sample <= -1040886;
 2994: sine_sample <= -1041079;
 2995: sine_sample <= -1041270;
 2996: sine_sample <= -1041458;
 2997: sine_sample <= -1041644;
 2998: sine_sample <= -1041828;
 2999: sine_sample <= -1042009;
 3000: sine_sample <= -1042187;
 3001: sine_sample <= -1042363;
 3002: sine_sample <= -1042537;
 3003: sine_sample <= -1042708;
 3004: sine_sample <= -1042877;
 3005: sine_sample <= -1043043;
 3006: sine_sample <= -1043207;
 3007: sine_sample <= -1043368;
 3008: sine_sample <= -1043527;
 3009: sine_sample <= -1043683;
 3010: sine_sample <= -1043837;
 3011: sine_sample <= -1043989;
 3012: sine_sample <= -1044138;
 3013: sine_sample <= -1044285;
 3014: sine_sample <= -1044429;
 3015: sine_sample <= -1044570;
 3016: sine_sample <= -1044710;
 3017: sine_sample <= -1044846;
 3018: sine_sample <= -1044981;
 3019: sine_sample <= -1045113;
 3020: sine_sample <= -1045242;
 3021: sine_sample <= -1045369;
 3022: sine_sample <= -1045493;
 3023: sine_sample <= -1045615;
 3024: sine_sample <= -1045735;
 3025: sine_sample <= -1045852;
 3026: sine_sample <= -1045967;
 3027: sine_sample <= -1046079;
 3028: sine_sample <= -1046189;
 3029: sine_sample <= -1046296;
 3030: sine_sample <= -1046401;
 3031: sine_sample <= -1046503;
 3032: sine_sample <= -1046603;
 3033: sine_sample <= -1046700;
 3034: sine_sample <= -1046795;
 3035: sine_sample <= -1046888;
 3036: sine_sample <= -1046978;
 3037: sine_sample <= -1047065;
 3038: sine_sample <= -1047150;
 3039: sine_sample <= -1047233;
 3040: sine_sample <= -1047313;
 3041: sine_sample <= -1047391;
 3042: sine_sample <= -1047466;
 3043: sine_sample <= -1047539;
 3044: sine_sample <= -1047609;
 3045: sine_sample <= -1047677;
 3046: sine_sample <= -1047742;
 3047: sine_sample <= -1047805;
 3048: sine_sample <= -1047866;
 3049: sine_sample <= -1047924;
 3050: sine_sample <= -1047979;
 3051: sine_sample <= -1048032;
 3052: sine_sample <= -1048083;
 3053: sine_sample <= -1048131;
 3054: sine_sample <= -1048176;
 3055: sine_sample <= -1048220;
 3056: sine_sample <= -1048260;
 3057: sine_sample <= -1048299;
 3058: sine_sample <= -1048334;
 3059: sine_sample <= -1048368;
 3060: sine_sample <= -1048398;
 3061: sine_sample <= -1048427;
 3062: sine_sample <= -1048453;
 3063: sine_sample <= -1048476;
 3064: sine_sample <= -1048497;
 3065: sine_sample <= -1048516;
 3066: sine_sample <= -1048532;
 3067: sine_sample <= -1048545;
 3068: sine_sample <= -1048556;
 3069: sine_sample <= -1048565;
 3070: sine_sample <= -1048571;
 3071: sine_sample <= -1048575;
 3072: sine_sample <= -1048576;
 3073: sine_sample <= -1048575;
 3074: sine_sample <= -1048571;
 3075: sine_sample <= -1048565;
 3076: sine_sample <= -1048556;
 3077: sine_sample <= -1048545;
 3078: sine_sample <= -1048532;
 3079: sine_sample <= -1048516;
 3080: sine_sample <= -1048497;
 3081: sine_sample <= -1048476;
 3082: sine_sample <= -1048453;
 3083: sine_sample <= -1048427;
 3084: sine_sample <= -1048398;
 3085: sine_sample <= -1048368;
 3086: sine_sample <= -1048334;
 3087: sine_sample <= -1048299;
 3088: sine_sample <= -1048260;
 3089: sine_sample <= -1048220;
 3090: sine_sample <= -1048176;
 3091: sine_sample <= -1048131;
 3092: sine_sample <= -1048083;
 3093: sine_sample <= -1048032;
 3094: sine_sample <= -1047979;
 3095: sine_sample <= -1047924;
 3096: sine_sample <= -1047866;
 3097: sine_sample <= -1047805;
 3098: sine_sample <= -1047742;
 3099: sine_sample <= -1047677;
 3100: sine_sample <= -1047609;
 3101: sine_sample <= -1047539;
 3102: sine_sample <= -1047466;
 3103: sine_sample <= -1047391;
 3104: sine_sample <= -1047313;
 3105: sine_sample <= -1047233;
 3106: sine_sample <= -1047150;
 3107: sine_sample <= -1047065;
 3108: sine_sample <= -1046978;
 3109: sine_sample <= -1046888;
 3110: sine_sample <= -1046795;
 3111: sine_sample <= -1046700;
 3112: sine_sample <= -1046603;
 3113: sine_sample <= -1046503;
 3114: sine_sample <= -1046401;
 3115: sine_sample <= -1046296;
 3116: sine_sample <= -1046189;
 3117: sine_sample <= -1046079;
 3118: sine_sample <= -1045967;
 3119: sine_sample <= -1045852;
 3120: sine_sample <= -1045735;
 3121: sine_sample <= -1045615;
 3122: sine_sample <= -1045493;
 3123: sine_sample <= -1045369;
 3124: sine_sample <= -1045242;
 3125: sine_sample <= -1045113;
 3126: sine_sample <= -1044981;
 3127: sine_sample <= -1044846;
 3128: sine_sample <= -1044710;
 3129: sine_sample <= -1044570;
 3130: sine_sample <= -1044429;
 3131: sine_sample <= -1044285;
 3132: sine_sample <= -1044138;
 3133: sine_sample <= -1043989;
 3134: sine_sample <= -1043837;
 3135: sine_sample <= -1043683;
 3136: sine_sample <= -1043527;
 3137: sine_sample <= -1043368;
 3138: sine_sample <= -1043207;
 3139: sine_sample <= -1043043;
 3140: sine_sample <= -1042877;
 3141: sine_sample <= -1042708;
 3142: sine_sample <= -1042537;
 3143: sine_sample <= -1042363;
 3144: sine_sample <= -1042187;
 3145: sine_sample <= -1042009;
 3146: sine_sample <= -1041828;
 3147: sine_sample <= -1041644;
 3148: sine_sample <= -1041458;
 3149: sine_sample <= -1041270;
 3150: sine_sample <= -1041079;
 3151: sine_sample <= -1040886;
 3152: sine_sample <= -1040690;
 3153: sine_sample <= -1040492;
 3154: sine_sample <= -1040292;
 3155: sine_sample <= -1040089;
 3156: sine_sample <= -1039883;
 3157: sine_sample <= -1039675;
 3158: sine_sample <= -1039465;
 3159: sine_sample <= -1039252;
 3160: sine_sample <= -1039037;
 3161: sine_sample <= -1038819;
 3162: sine_sample <= -1038599;
 3163: sine_sample <= -1038376;
 3164: sine_sample <= -1038151;
 3165: sine_sample <= -1037924;
 3166: sine_sample <= -1037694;
 3167: sine_sample <= -1037462;
 3168: sine_sample <= -1037227;
 3169: sine_sample <= -1036990;
 3170: sine_sample <= -1036750;
 3171: sine_sample <= -1036508;
 3172: sine_sample <= -1036263;
 3173: sine_sample <= -1036016;
 3174: sine_sample <= -1035767;
 3175: sine_sample <= -1035515;
 3176: sine_sample <= -1035261;
 3177: sine_sample <= -1035004;
 3178: sine_sample <= -1034745;
 3179: sine_sample <= -1034483;
 3180: sine_sample <= -1034219;
 3181: sine_sample <= -1033953;
 3182: sine_sample <= -1033684;
 3183: sine_sample <= -1033412;
 3184: sine_sample <= -1033139;
 3185: sine_sample <= -1032862;
 3186: sine_sample <= -1032584;
 3187: sine_sample <= -1032303;
 3188: sine_sample <= -1032019;
 3189: sine_sample <= -1031733;
 3190: sine_sample <= -1031445;
 3191: sine_sample <= -1031154;
 3192: sine_sample <= -1030861;
 3193: sine_sample <= -1030565;
 3194: sine_sample <= -1030267;
 3195: sine_sample <= -1029967;
 3196: sine_sample <= -1029664;
 3197: sine_sample <= -1029359;
 3198: sine_sample <= -1029051;
 3199: sine_sample <= -1028741;
 3200: sine_sample <= -1028428;
 3201: sine_sample <= -1028113;
 3202: sine_sample <= -1027796;
 3203: sine_sample <= -1027476;
 3204: sine_sample <= -1027153;
 3205: sine_sample <= -1026829;
 3206: sine_sample <= -1026502;
 3207: sine_sample <= -1026172;
 3208: sine_sample <= -1025840;
 3209: sine_sample <= -1025506;
 3210: sine_sample <= -1025169;
 3211: sine_sample <= -1024830;
 3212: sine_sample <= -1024488;
 3213: sine_sample <= -1024144;
 3214: sine_sample <= -1023798;
 3215: sine_sample <= -1023449;
 3216: sine_sample <= -1023098;
 3217: sine_sample <= -1022744;
 3218: sine_sample <= -1022388;
 3219: sine_sample <= -1022030;
 3220: sine_sample <= -1021669;
 3221: sine_sample <= -1021306;
 3222: sine_sample <= -1020940;
 3223: sine_sample <= -1020572;
 3224: sine_sample <= -1020202;
 3225: sine_sample <= -1019829;
 3226: sine_sample <= -1019453;
 3227: sine_sample <= -1019076;
 3228: sine_sample <= -1018696;
 3229: sine_sample <= -1018313;
 3230: sine_sample <= -1017928;
 3231: sine_sample <= -1017541;
 3232: sine_sample <= -1017152;
 3233: sine_sample <= -1016760;
 3234: sine_sample <= -1016365;
 3235: sine_sample <= -1015968;
 3236: sine_sample <= -1015569;
 3237: sine_sample <= -1015168;
 3238: sine_sample <= -1014764;
 3239: sine_sample <= -1014357;
 3240: sine_sample <= -1013948;
 3241: sine_sample <= -1013537;
 3242: sine_sample <= -1013124;
 3243: sine_sample <= -1012708;
 3244: sine_sample <= -1012290;
 3245: sine_sample <= -1011869;
 3246: sine_sample <= -1011446;
 3247: sine_sample <= -1011020;
 3248: sine_sample <= -1010593;
 3249: sine_sample <= -1010162;
 3250: sine_sample <= -1009730;
 3251: sine_sample <= -1009295;
 3252: sine_sample <= -1008858;
 3253: sine_sample <= -1008418;
 3254: sine_sample <= -1007976;
 3255: sine_sample <= -1007531;
 3256: sine_sample <= -1007085;
 3257: sine_sample <= -1006635;
 3258: sine_sample <= -1006184;
 3259: sine_sample <= -1005730;
 3260: sine_sample <= -1005274;
 3261: sine_sample <= -1004815;
 3262: sine_sample <= -1004354;
 3263: sine_sample <= -1003891;
 3264: sine_sample <= -1003425;
 3265: sine_sample <= -1002957;
 3266: sine_sample <= -1002486;
 3267: sine_sample <= -1002013;
 3268: sine_sample <= -1001538;
 3269: sine_sample <= -1001061;
 3270: sine_sample <= -1000581;
 3271: sine_sample <= -1000099;
 3272: sine_sample <= -999614;
 3273: sine_sample <= -999127;
 3274: sine_sample <= -998638;
 3275: sine_sample <= -998146;
 3276: sine_sample <= -997652;
 3277: sine_sample <= -997156;
 3278: sine_sample <= -996657;
 3279: sine_sample <= -996156;
 3280: sine_sample <= -995653;
 3281: sine_sample <= -995147;
 3282: sine_sample <= -994639;
 3283: sine_sample <= -994128;
 3284: sine_sample <= -993616;
 3285: sine_sample <= -993101;
 3286: sine_sample <= -992583;
 3287: sine_sample <= -992063;
 3288: sine_sample <= -991541;
 3289: sine_sample <= -991017;
 3290: sine_sample <= -990490;
 3291: sine_sample <= -989961;
 3292: sine_sample <= -989430;
 3293: sine_sample <= -988896;
 3294: sine_sample <= -988360;
 3295: sine_sample <= -987821;
 3296: sine_sample <= -987281;
 3297: sine_sample <= -986738;
 3298: sine_sample <= -986192;
 3299: sine_sample <= -985645;
 3300: sine_sample <= -985095;
 3301: sine_sample <= -984542;
 3302: sine_sample <= -983988;
 3303: sine_sample <= -983431;
 3304: sine_sample <= -982871;
 3305: sine_sample <= -982310;
 3306: sine_sample <= -981746;
 3307: sine_sample <= -981180;
 3308: sine_sample <= -980611;
 3309: sine_sample <= -980040;
 3310: sine_sample <= -979467;
 3311: sine_sample <= -978892;
 3312: sine_sample <= -978314;
 3313: sine_sample <= -977734;
 3314: sine_sample <= -977152;
 3315: sine_sample <= -976567;
 3316: sine_sample <= -975980;
 3317: sine_sample <= -975391;
 3318: sine_sample <= -974799;
 3319: sine_sample <= -974205;
 3320: sine_sample <= -973609;
 3321: sine_sample <= -973011;
 3322: sine_sample <= -972410;
 3323: sine_sample <= -971807;
 3324: sine_sample <= -971202;
 3325: sine_sample <= -970594;
 3326: sine_sample <= -969985;
 3327: sine_sample <= -969372;
 3328: sine_sample <= -968758;
 3329: sine_sample <= -968141;
 3330: sine_sample <= -967522;
 3331: sine_sample <= -966901;
 3332: sine_sample <= -966278;
 3333: sine_sample <= -965652;
 3334: sine_sample <= -965024;
 3335: sine_sample <= -964393;
 3336: sine_sample <= -963761;
 3337: sine_sample <= -963126;
 3338: sine_sample <= -962489;
 3339: sine_sample <= -961849;
 3340: sine_sample <= -961208;
 3341: sine_sample <= -960564;
 3342: sine_sample <= -959918;
 3343: sine_sample <= -959269;
 3344: sine_sample <= -958619;
 3345: sine_sample <= -957966;
 3346: sine_sample <= -957310;
 3347: sine_sample <= -956653;
 3348: sine_sample <= -955993;
 3349: sine_sample <= -955331;
 3350: sine_sample <= -954667;
 3351: sine_sample <= -954001;
 3352: sine_sample <= -953332;
 3353: sine_sample <= -952661;
 3354: sine_sample <= -951988;
 3355: sine_sample <= -951312;
 3356: sine_sample <= -950635;
 3357: sine_sample <= -949955;
 3358: sine_sample <= -949273;
 3359: sine_sample <= -948588;
 3360: sine_sample <= -947902;
 3361: sine_sample <= -947213;
 3362: sine_sample <= -946522;
 3363: sine_sample <= -945828;
 3364: sine_sample <= -945133;
 3365: sine_sample <= -944435;
 3366: sine_sample <= -943735;
 3367: sine_sample <= -943033;
 3368: sine_sample <= -942329;
 3369: sine_sample <= -941622;
 3370: sine_sample <= -940913;
 3371: sine_sample <= -940202;
 3372: sine_sample <= -939489;
 3373: sine_sample <= -938773;
 3374: sine_sample <= -938056;
 3375: sine_sample <= -937336;
 3376: sine_sample <= -936614;
 3377: sine_sample <= -935889;
 3378: sine_sample <= -935163;
 3379: sine_sample <= -934434;
 3380: sine_sample <= -933703;
 3381: sine_sample <= -932970;
 3382: sine_sample <= -932235;
 3383: sine_sample <= -931497;
 3384: sine_sample <= -930758;
 3385: sine_sample <= -930016;
 3386: sine_sample <= -929272;
 3387: sine_sample <= -928526;
 3388: sine_sample <= -927777;
 3389: sine_sample <= -927027;
 3390: sine_sample <= -926274;
 3391: sine_sample <= -925519;
 3392: sine_sample <= -924762;
 3393: sine_sample <= -924002;
 3394: sine_sample <= -923241;
 3395: sine_sample <= -922477;
 3396: sine_sample <= -921711;
 3397: sine_sample <= -920943;
 3398: sine_sample <= -920173;
 3399: sine_sample <= -919401;
 3400: sine_sample <= -918626;
 3401: sine_sample <= -917850;
 3402: sine_sample <= -917071;
 3403: sine_sample <= -916290;
 3404: sine_sample <= -915507;
 3405: sine_sample <= -914721;
 3406: sine_sample <= -913934;
 3407: sine_sample <= -913144;
 3408: sine_sample <= -912352;
 3409: sine_sample <= -911559;
 3410: sine_sample <= -910763;
 3411: sine_sample <= -909964;
 3412: sine_sample <= -909164;
 3413: sine_sample <= -908362;
 3414: sine_sample <= -907557;
 3415: sine_sample <= -906750;
 3416: sine_sample <= -905941;
 3417: sine_sample <= -905130;
 3418: sine_sample <= -904317;
 3419: sine_sample <= -903502;
 3420: sine_sample <= -902685;
 3421: sine_sample <= -901865;
 3422: sine_sample <= -901043;
 3423: sine_sample <= -900220;
 3424: sine_sample <= -899394;
 3425: sine_sample <= -898566;
 3426: sine_sample <= -897736;
 3427: sine_sample <= -896903;
 3428: sine_sample <= -896069;
 3429: sine_sample <= -895233;
 3430: sine_sample <= -894394;
 3431: sine_sample <= -893553;
 3432: sine_sample <= -892711;
 3433: sine_sample <= -891866;
 3434: sine_sample <= -891019;
 3435: sine_sample <= -890170;
 3436: sine_sample <= -889319;
 3437: sine_sample <= -888466;
 3438: sine_sample <= -887610;
 3439: sine_sample <= -886753;
 3440: sine_sample <= -885893;
 3441: sine_sample <= -885032;
 3442: sine_sample <= -884168;
 3443: sine_sample <= -883302;
 3444: sine_sample <= -882434;
 3445: sine_sample <= -881565;
 3446: sine_sample <= -880693;
 3447: sine_sample <= -879819;
 3448: sine_sample <= -878942;
 3449: sine_sample <= -878064;
 3450: sine_sample <= -877184;
 3451: sine_sample <= -876302;
 3452: sine_sample <= -875417;
 3453: sine_sample <= -874531;
 3454: sine_sample <= -873642;
 3455: sine_sample <= -872752;
 3456: sine_sample <= -871859;
 3457: sine_sample <= -870965;
 3458: sine_sample <= -870068;
 3459: sine_sample <= -869169;
 3460: sine_sample <= -868268;
 3461: sine_sample <= -867365;
 3462: sine_sample <= -866461;
 3463: sine_sample <= -865554;
 3464: sine_sample <= -864645;
 3465: sine_sample <= -863734;
 3466: sine_sample <= -862821;
 3467: sine_sample <= -861906;
 3468: sine_sample <= -860989;
 3469: sine_sample <= -860069;
 3470: sine_sample <= -859148;
 3471: sine_sample <= -858225;
 3472: sine_sample <= -857300;
 3473: sine_sample <= -856373;
 3474: sine_sample <= -855444;
 3475: sine_sample <= -854512;
 3476: sine_sample <= -853579;
 3477: sine_sample <= -852644;
 3478: sine_sample <= -851707;
 3479: sine_sample <= -850767;
 3480: sine_sample <= -849826;
 3481: sine_sample <= -848883;
 3482: sine_sample <= -847938;
 3483: sine_sample <= -846990;
 3484: sine_sample <= -846041;
 3485: sine_sample <= -845090;
 3486: sine_sample <= -844137;
 3487: sine_sample <= -843181;
 3488: sine_sample <= -842224;
 3489: sine_sample <= -841265;
 3490: sine_sample <= -840304;
 3491: sine_sample <= -839341;
 3492: sine_sample <= -838376;
 3493: sine_sample <= -837409;
 3494: sine_sample <= -836440;
 3495: sine_sample <= -835469;
 3496: sine_sample <= -834496;
 3497: sine_sample <= -833521;
 3498: sine_sample <= -832544;
 3499: sine_sample <= -831565;
 3500: sine_sample <= -830584;
 3501: sine_sample <= -829601;
 3502: sine_sample <= -828617;
 3503: sine_sample <= -827630;
 3504: sine_sample <= -826641;
 3505: sine_sample <= -825651;
 3506: sine_sample <= -824658;
 3507: sine_sample <= -823664;
 3508: sine_sample <= -822667;
 3509: sine_sample <= -821669;
 3510: sine_sample <= -820669;
 3511: sine_sample <= -819667;
 3512: sine_sample <= -818662;
 3513: sine_sample <= -817656;
 3514: sine_sample <= -816648;
 3515: sine_sample <= -815639;
 3516: sine_sample <= -814627;
 3517: sine_sample <= -813613;
 3518: sine_sample <= -812597;
 3519: sine_sample <= -811580;
 3520: sine_sample <= -810560;
 3521: sine_sample <= -809539;
 3522: sine_sample <= -808516;
 3523: sine_sample <= -807491;
 3524: sine_sample <= -806463;
 3525: sine_sample <= -805434;
 3526: sine_sample <= -804404;
 3527: sine_sample <= -803371;
 3528: sine_sample <= -802336;
 3529: sine_sample <= -801300;
 3530: sine_sample <= -800261;
 3531: sine_sample <= -799221;
 3532: sine_sample <= -798179;
 3533: sine_sample <= -797135;
 3534: sine_sample <= -796089;
 3535: sine_sample <= -795041;
 3536: sine_sample <= -793991;
 3537: sine_sample <= -792940;
 3538: sine_sample <= -791886;
 3539: sine_sample <= -790831;
 3540: sine_sample <= -789774;
 3541: sine_sample <= -788715;
 3542: sine_sample <= -787654;
 3543: sine_sample <= -786591;
 3544: sine_sample <= -785527;
 3545: sine_sample <= -784460;
 3546: sine_sample <= -783392;
 3547: sine_sample <= -782322;
 3548: sine_sample <= -781250;
 3549: sine_sample <= -780176;
 3550: sine_sample <= -779100;
 3551: sine_sample <= -778023;
 3552: sine_sample <= -776944;
 3553: sine_sample <= -775863;
 3554: sine_sample <= -774780;
 3555: sine_sample <= -773695;
 3556: sine_sample <= -772608;
 3557: sine_sample <= -771520;
 3558: sine_sample <= -770430;
 3559: sine_sample <= -769338;
 3560: sine_sample <= -768244;
 3561: sine_sample <= -767148;
 3562: sine_sample <= -766051;
 3563: sine_sample <= -764951;
 3564: sine_sample <= -763850;
 3565: sine_sample <= -762748;
 3566: sine_sample <= -761643;
 3567: sine_sample <= -760536;
 3568: sine_sample <= -759428;
 3569: sine_sample <= -758318;
 3570: sine_sample <= -757206;
 3571: sine_sample <= -756093;
 3572: sine_sample <= -754977;
 3573: sine_sample <= -753860;
 3574: sine_sample <= -752741;
 3575: sine_sample <= -751621;
 3576: sine_sample <= -750498;
 3577: sine_sample <= -749374;
 3578: sine_sample <= -748248;
 3579: sine_sample <= -747120;
 3580: sine_sample <= -745991;
 3581: sine_sample <= -744860;
 3582: sine_sample <= -743727;
 3583: sine_sample <= -742592;
 3584: sine_sample <= -741455;
 3585: sine_sample <= -740317;
 3586: sine_sample <= -739177;
 3587: sine_sample <= -738035;
 3588: sine_sample <= -736892;
 3589: sine_sample <= -735747;
 3590: sine_sample <= -734600;
 3591: sine_sample <= -733451;
 3592: sine_sample <= -732301;
 3593: sine_sample <= -731149;
 3594: sine_sample <= -729995;
 3595: sine_sample <= -728839;
 3596: sine_sample <= -727682;
 3597: sine_sample <= -726523;
 3598: sine_sample <= -725362;
 3599: sine_sample <= -724200;
 3600: sine_sample <= -723036;
 3601: sine_sample <= -721870;
 3602: sine_sample <= -720702;
 3603: sine_sample <= -719533;
 3604: sine_sample <= -718362;
 3605: sine_sample <= -717190;
 3606: sine_sample <= -716016;
 3607: sine_sample <= -714840;
 3608: sine_sample <= -713662;
 3609: sine_sample <= -712483;
 3610: sine_sample <= -711302;
 3611: sine_sample <= -710119;
 3612: sine_sample <= -708935;
 3613: sine_sample <= -707749;
 3614: sine_sample <= -706561;
 3615: sine_sample <= -705372;
 3616: sine_sample <= -704181;
 3617: sine_sample <= -702988;
 3618: sine_sample <= -701794;
 3619: sine_sample <= -700598;
 3620: sine_sample <= -699400;
 3621: sine_sample <= -698201;
 3622: sine_sample <= -697000;
 3623: sine_sample <= -695798;
 3624: sine_sample <= -694593;
 3625: sine_sample <= -693388;
 3626: sine_sample <= -692180;
 3627: sine_sample <= -690971;
 3628: sine_sample <= -689760;
 3629: sine_sample <= -688548;
 3630: sine_sample <= -687334;
 3631: sine_sample <= -686119;
 3632: sine_sample <= -684901;
 3633: sine_sample <= -683683;
 3634: sine_sample <= -682462;
 3635: sine_sample <= -681240;
 3636: sine_sample <= -680017;
 3637: sine_sample <= -678792;
 3638: sine_sample <= -677565;
 3639: sine_sample <= -676336;
 3640: sine_sample <= -675106;
 3641: sine_sample <= -673875;
 3642: sine_sample <= -672642;
 3643: sine_sample <= -671407;
 3644: sine_sample <= -670171;
 3645: sine_sample <= -668933;
 3646: sine_sample <= -667693;
 3647: sine_sample <= -666452;
 3648: sine_sample <= -665210;
 3649: sine_sample <= -663966;
 3650: sine_sample <= -662720;
 3651: sine_sample <= -661473;
 3652: sine_sample <= -660224;
 3653: sine_sample <= -658973;
 3654: sine_sample <= -657721;
 3655: sine_sample <= -656468;
 3656: sine_sample <= -655213;
 3657: sine_sample <= -653956;
 3658: sine_sample <= -652698;
 3659: sine_sample <= -651438;
 3660: sine_sample <= -650177;
 3661: sine_sample <= -648915;
 3662: sine_sample <= -647650;
 3663: sine_sample <= -646384;
 3664: sine_sample <= -645117;
 3665: sine_sample <= -643848;
 3666: sine_sample <= -642578;
 3667: sine_sample <= -641306;
 3668: sine_sample <= -640033;
 3669: sine_sample <= -638758;
 3670: sine_sample <= -637482;
 3671: sine_sample <= -636204;
 3672: sine_sample <= -634924;
 3673: sine_sample <= -633644;
 3674: sine_sample <= -632361;
 3675: sine_sample <= -631077;
 3676: sine_sample <= -629792;
 3677: sine_sample <= -628505;
 3678: sine_sample <= -627217;
 3679: sine_sample <= -625927;
 3680: sine_sample <= -624636;
 3681: sine_sample <= -623343;
 3682: sine_sample <= -622049;
 3683: sine_sample <= -620754;
 3684: sine_sample <= -619457;
 3685: sine_sample <= -618158;
 3686: sine_sample <= -616858;
 3687: sine_sample <= -615557;
 3688: sine_sample <= -614254;
 3689: sine_sample <= -612949;
 3690: sine_sample <= -611644;
 3691: sine_sample <= -610336;
 3692: sine_sample <= -609028;
 3693: sine_sample <= -607718;
 3694: sine_sample <= -606406;
 3695: sine_sample <= -605093;
 3696: sine_sample <= -603779;
 3697: sine_sample <= -602463;
 3698: sine_sample <= -601146;
 3699: sine_sample <= -599827;
 3700: sine_sample <= -598507;
 3701: sine_sample <= -597186;
 3702: sine_sample <= -595863;
 3703: sine_sample <= -594539;
 3704: sine_sample <= -593213;
 3705: sine_sample <= -591886;
 3706: sine_sample <= -590557;
 3707: sine_sample <= -589228;
 3708: sine_sample <= -587896;
 3709: sine_sample <= -586564;
 3710: sine_sample <= -585230;
 3711: sine_sample <= -583894;
 3712: sine_sample <= -582558;
 3713: sine_sample <= -581220;
 3714: sine_sample <= -579880;
 3715: sine_sample <= -578539;
 3716: sine_sample <= -577197;
 3717: sine_sample <= -575854;
 3718: sine_sample <= -574509;
 3719: sine_sample <= -573162;
 3720: sine_sample <= -571815;
 3721: sine_sample <= -570466;
 3722: sine_sample <= -569116;
 3723: sine_sample <= -567764;
 3724: sine_sample <= -566411;
 3725: sine_sample <= -565057;
 3726: sine_sample <= -563701;
 3727: sine_sample <= -562344;
 3728: sine_sample <= -560986;
 3729: sine_sample <= -559626;
 3730: sine_sample <= -558265;
 3731: sine_sample <= -556903;
 3732: sine_sample <= -555539;
 3733: sine_sample <= -554175;
 3734: sine_sample <= -552808;
 3735: sine_sample <= -551441;
 3736: sine_sample <= -550072;
 3737: sine_sample <= -548702;
 3738: sine_sample <= -547331;
 3739: sine_sample <= -545958;
 3740: sine_sample <= -544584;
 3741: sine_sample <= -543209;
 3742: sine_sample <= -541833;
 3743: sine_sample <= -540455;
 3744: sine_sample <= -539076;
 3745: sine_sample <= -537696;
 3746: sine_sample <= -536314;
 3747: sine_sample <= -534931;
 3748: sine_sample <= -533547;
 3749: sine_sample <= -532162;
 3750: sine_sample <= -530775;
 3751: sine_sample <= -529387;
 3752: sine_sample <= -527998;
 3753: sine_sample <= -526608;
 3754: sine_sample <= -525217;
 3755: sine_sample <= -523824;
 3756: sine_sample <= -522430;
 3757: sine_sample <= -521034;
 3758: sine_sample <= -519638;
 3759: sine_sample <= -518240;
 3760: sine_sample <= -516841;
 3761: sine_sample <= -515441;
 3762: sine_sample <= -514040;
 3763: sine_sample <= -512637;
 3764: sine_sample <= -511234;
 3765: sine_sample <= -509829;
 3766: sine_sample <= -508422;
 3767: sine_sample <= -507015;
 3768: sine_sample <= -505606;
 3769: sine_sample <= -504197;
 3770: sine_sample <= -502786;
 3771: sine_sample <= -501374;
 3772: sine_sample <= -499960;
 3773: sine_sample <= -498546;
 3774: sine_sample <= -497130;
 3775: sine_sample <= -495713;
 3776: sine_sample <= -494295;
 3777: sine_sample <= -492876;
 3778: sine_sample <= -491456;
 3779: sine_sample <= -490035;
 3780: sine_sample <= -488612;
 3781: sine_sample <= -487188;
 3782: sine_sample <= -485763;
 3783: sine_sample <= -484337;
 3784: sine_sample <= -482910;
 3785: sine_sample <= -481482;
 3786: sine_sample <= -480052;
 3787: sine_sample <= -478622;
 3788: sine_sample <= -477190;
 3789: sine_sample <= -475757;
 3790: sine_sample <= -474323;
 3791: sine_sample <= -472888;
 3792: sine_sample <= -471452;
 3793: sine_sample <= -470014;
 3794: sine_sample <= -468576;
 3795: sine_sample <= -467137;
 3796: sine_sample <= -465696;
 3797: sine_sample <= -464254;
 3798: sine_sample <= -462811;
 3799: sine_sample <= -461368;
 3800: sine_sample <= -459923;
 3801: sine_sample <= -458477;
 3802: sine_sample <= -457029;
 3803: sine_sample <= -455581;
 3804: sine_sample <= -454132;
 3805: sine_sample <= -452682;
 3806: sine_sample <= -451230;
 3807: sine_sample <= -449778;
 3808: sine_sample <= -448324;
 3809: sine_sample <= -446870;
 3810: sine_sample <= -445414;
 3811: sine_sample <= -443957;
 3812: sine_sample <= -442499;
 3813: sine_sample <= -441041;
 3814: sine_sample <= -439581;
 3815: sine_sample <= -438120;
 3816: sine_sample <= -436658;
 3817: sine_sample <= -435195;
 3818: sine_sample <= -433731;
 3819: sine_sample <= -432266;
 3820: sine_sample <= -430800;
 3821: sine_sample <= -429333;
 3822: sine_sample <= -427865;
 3823: sine_sample <= -426396;
 3824: sine_sample <= -424926;
 3825: sine_sample <= -423455;
 3826: sine_sample <= -421983;
 3827: sine_sample <= -420510;
 3828: sine_sample <= -419036;
 3829: sine_sample <= -417562;
 3830: sine_sample <= -416086;
 3831: sine_sample <= -414609;
 3832: sine_sample <= -413131;
 3833: sine_sample <= -411652;
 3834: sine_sample <= -410172;
 3835: sine_sample <= -408691;
 3836: sine_sample <= -407209;
 3837: sine_sample <= -405727;
 3838: sine_sample <= -404243;
 3839: sine_sample <= -402758;
 3840: sine_sample <= -401273;
 3841: sine_sample <= -399786;
 3842: sine_sample <= -398299;
 3843: sine_sample <= -396810;
 3844: sine_sample <= -395321;
 3845: sine_sample <= -393831;
 3846: sine_sample <= -392340;
 3847: sine_sample <= -390847;
 3848: sine_sample <= -389354;
 3849: sine_sample <= -387860;
 3850: sine_sample <= -386366;
 3851: sine_sample <= -384870;
 3852: sine_sample <= -383373;
 3853: sine_sample <= -381876;
 3854: sine_sample <= -380377;
 3855: sine_sample <= -378878;
 3856: sine_sample <= -377377;
 3857: sine_sample <= -375876;
 3858: sine_sample <= -374374;
 3859: sine_sample <= -372871;
 3860: sine_sample <= -371367;
 3861: sine_sample <= -369863;
 3862: sine_sample <= -368357;
 3863: sine_sample <= -366851;
 3864: sine_sample <= -365344;
 3865: sine_sample <= -363835;
 3866: sine_sample <= -362326;
 3867: sine_sample <= -360817;
 3868: sine_sample <= -359306;
 3869: sine_sample <= -357794;
 3870: sine_sample <= -356282;
 3871: sine_sample <= -354769;
 3872: sine_sample <= -353255;
 3873: sine_sample <= -351740;
 3874: sine_sample <= -350224;
 3875: sine_sample <= -348708;
 3876: sine_sample <= -347190;
 3877: sine_sample <= -345672;
 3878: sine_sample <= -344153;
 3879: sine_sample <= -342633;
 3880: sine_sample <= -341113;
 3881: sine_sample <= -339591;
 3882: sine_sample <= -338069;
 3883: sine_sample <= -336546;
 3884: sine_sample <= -335022;
 3885: sine_sample <= -333498;
 3886: sine_sample <= -331972;
 3887: sine_sample <= -330446;
 3888: sine_sample <= -328919;
 3889: sine_sample <= -327392;
 3890: sine_sample <= -325863;
 3891: sine_sample <= -324334;
 3892: sine_sample <= -322804;
 3893: sine_sample <= -321273;
 3894: sine_sample <= -319742;
 3895: sine_sample <= -318209;
 3896: sine_sample <= -316676;
 3897: sine_sample <= -315143;
 3898: sine_sample <= -313608;
 3899: sine_sample <= -312073;
 3900: sine_sample <= -310537;
 3901: sine_sample <= -309000;
 3902: sine_sample <= -307463;
 3903: sine_sample <= -305925;
 3904: sine_sample <= -304386;
 3905: sine_sample <= -302846;
 3906: sine_sample <= -301306;
 3907: sine_sample <= -299765;
 3908: sine_sample <= -298223;
 3909: sine_sample <= -296681;
 3910: sine_sample <= -295138;
 3911: sine_sample <= -293594;
 3912: sine_sample <= -292049;
 3913: sine_sample <= -290504;
 3914: sine_sample <= -288958;
 3915: sine_sample <= -287412;
 3916: sine_sample <= -285864;
 3917: sine_sample <= -284316;
 3918: sine_sample <= -282768;
 3919: sine_sample <= -281219;
 3920: sine_sample <= -279669;
 3921: sine_sample <= -278118;
 3922: sine_sample <= -276567;
 3923: sine_sample <= -275015;
 3924: sine_sample <= -273463;
 3925: sine_sample <= -271909;
 3926: sine_sample <= -270356;
 3927: sine_sample <= -268801;
 3928: sine_sample <= -267246;
 3929: sine_sample <= -265690;
 3930: sine_sample <= -264134;
 3931: sine_sample <= -262577;
 3932: sine_sample <= -261020;
 3933: sine_sample <= -259461;
 3934: sine_sample <= -257903;
 3935: sine_sample <= -256343;
 3936: sine_sample <= -254783;
 3937: sine_sample <= -253223;
 3938: sine_sample <= -251662;
 3939: sine_sample <= -250100;
 3940: sine_sample <= -248537;
 3941: sine_sample <= -246974;
 3942: sine_sample <= -245411;
 3943: sine_sample <= -243847;
 3944: sine_sample <= -242282;
 3945: sine_sample <= -240717;
 3946: sine_sample <= -239151;
 3947: sine_sample <= -237585;
 3948: sine_sample <= -236018;
 3949: sine_sample <= -234450;
 3950: sine_sample <= -232882;
 3951: sine_sample <= -231314;
 3952: sine_sample <= -229744;
 3953: sine_sample <= -228175;
 3954: sine_sample <= -226605;
 3955: sine_sample <= -225034;
 3956: sine_sample <= -223462;
 3957: sine_sample <= -221891;
 3958: sine_sample <= -220318;
 3959: sine_sample <= -218746;
 3960: sine_sample <= -217172;
 3961: sine_sample <= -215598;
 3962: sine_sample <= -214024;
 3963: sine_sample <= -212449;
 3964: sine_sample <= -210874;
 3965: sine_sample <= -209298;
 3966: sine_sample <= -207721;
 3967: sine_sample <= -206145;
 3968: sine_sample <= -204567;
 3969: sine_sample <= -202989;
 3970: sine_sample <= -201411;
 3971: sine_sample <= -199832;
 3972: sine_sample <= -198253;
 3973: sine_sample <= -196673;
 3974: sine_sample <= -195093;
 3975: sine_sample <= -193512;
 3976: sine_sample <= -191931;
 3977: sine_sample <= -190350;
 3978: sine_sample <= -188768;
 3979: sine_sample <= -187185;
 3980: sine_sample <= -185603;
 3981: sine_sample <= -184019;
 3982: sine_sample <= -182435;
 3983: sine_sample <= -180851;
 3984: sine_sample <= -179267;
 3985: sine_sample <= -177682;
 3986: sine_sample <= -176096;
 3987: sine_sample <= -174510;
 3988: sine_sample <= -172924;
 3989: sine_sample <= -171337;
 3990: sine_sample <= -169750;
 3991: sine_sample <= -168163;
 3992: sine_sample <= -166575;
 3993: sine_sample <= -164987;
 3994: sine_sample <= -163398;
 3995: sine_sample <= -161809;
 3996: sine_sample <= -160220;
 3997: sine_sample <= -158630;
 3998: sine_sample <= -157040;
 3999: sine_sample <= -155449;
 4000: sine_sample <= -153858;
 4001: sine_sample <= -152267;
 4002: sine_sample <= -150675;
 4003: sine_sample <= -149083;
 4004: sine_sample <= -147491;
 4005: sine_sample <= -145898;
 4006: sine_sample <= -144305;
 4007: sine_sample <= -142712;
 4008: sine_sample <= -141118;
 4009: sine_sample <= -139524;
 4010: sine_sample <= -137930;
 4011: sine_sample <= -136335;
 4012: sine_sample <= -134740;
 4013: sine_sample <= -133145;
 4014: sine_sample <= -131549;
 4015: sine_sample <= -129953;
 4016: sine_sample <= -128357;
 4017: sine_sample <= -126760;
 4018: sine_sample <= -125164;
 4019: sine_sample <= -123566;
 4020: sine_sample <= -121969;
 4021: sine_sample <= -120371;
 4022: sine_sample <= -118773;
 4023: sine_sample <= -117175;
 4024: sine_sample <= -115576;
 4025: sine_sample <= -113978;
 4026: sine_sample <= -112379;
 4027: sine_sample <= -110779;
 4028: sine_sample <= -109180;
 4029: sine_sample <= -107580;
 4030: sine_sample <= -105980;
 4031: sine_sample <= -104379;
 4032: sine_sample <= -102779;
 4033: sine_sample <= -101178;
 4034: sine_sample <= -99577;
 4035: sine_sample <= -97975;
 4036: sine_sample <= -96374;
 4037: sine_sample <= -94772;
 4038: sine_sample <= -93170;
 4039: sine_sample <= -91568;
 4040: sine_sample <= -89965;
 4041: sine_sample <= -88362;
 4042: sine_sample <= -86760;
 4043: sine_sample <= -85156;
 4044: sine_sample <= -83553;
 4045: sine_sample <= -81950;
 4046: sine_sample <= -80346;
 4047: sine_sample <= -78742;
 4048: sine_sample <= -77138;
 4049: sine_sample <= -75534;
 4050: sine_sample <= -73930;
 4051: sine_sample <= -72325;
 4052: sine_sample <= -70720;
 4053: sine_sample <= -69115;
 4054: sine_sample <= -67510;
 4055: sine_sample <= -65905;
 4056: sine_sample <= -64300;
 4057: sine_sample <= -62694;
 4058: sine_sample <= -61088;
 4059: sine_sample <= -59483;
 4060: sine_sample <= -57877;
 4061: sine_sample <= -56270;
 4062: sine_sample <= -54664;
 4063: sine_sample <= -53058;
 4064: sine_sample <= -51451;
 4065: sine_sample <= -49845;
 4066: sine_sample <= -48238;
 4067: sine_sample <= -46631;
 4068: sine_sample <= -45024;
 4069: sine_sample <= -43417;
 4070: sine_sample <= -41810;
 4071: sine_sample <= -40203;
 4072: sine_sample <= -38595;
 4073: sine_sample <= -36988;
 4074: sine_sample <= -35380;
 4075: sine_sample <= -33773;
 4076: sine_sample <= -32165;
 4077: sine_sample <= -30557;
 4078: sine_sample <= -28949;
 4079: sine_sample <= -27341;
 4080: sine_sample <= -25733;
 4081: sine_sample <= -24125;
 4082: sine_sample <= -22517;
 4083: sine_sample <= -20909;
 4084: sine_sample <= -19301;
 4085: sine_sample <= -17693;
 4086: sine_sample <= -16084;
 4087: sine_sample <= -14476;
 4088: sine_sample <= -12868;
 4089: sine_sample <= -11259;
 4090: sine_sample <= -9651;
 4091: sine_sample <= -8043;
 4092: sine_sample <= -6434;
 4093: sine_sample <= -4826;
 4094: sine_sample <= -3217;
 4095: sine_sample <= -1609;
 default: sine_sample <= 24'b0;
 endcase
 end

assign dout = sine_sample;

 endmodule 